library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
entity project_tb is
end project_tb;
architecture projecttb of project_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;
type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (
			0 => std_logic_vector(to_unsigned(16, 8)),
			1 => std_logic_vector(to_unsigned(71, 8)),
			2 => std_logic_vector(to_unsigned(14, 8)),
			3 => std_logic_vector(to_unsigned(207, 8)),
			4 => std_logic_vector(to_unsigned(248, 8)),
			5 => std_logic_vector(to_unsigned(169, 8)),
			6 => std_logic_vector(to_unsigned(34, 8)),
			7 => std_logic_vector(to_unsigned(19, 8)),
			8 => std_logic_vector(to_unsigned(108, 8)),
			9 => std_logic_vector(to_unsigned(54, 8)),
			10 => std_logic_vector(to_unsigned(36, 8)),
			11 => std_logic_vector(to_unsigned(162, 8)),
			12 => std_logic_vector(to_unsigned(190, 8)),
			13 => std_logic_vector(to_unsigned(105, 8)),
			14 => std_logic_vector(to_unsigned(202, 8)),
			15 => std_logic_vector(to_unsigned(160, 8)),
			16 => std_logic_vector(to_unsigned(215, 8)),
			17 => std_logic_vector(to_unsigned(158, 8)),
			18 => std_logic_vector(to_unsigned(203, 8)),
			19 => std_logic_vector(to_unsigned(78, 8)),
			20 => std_logic_vector(to_unsigned(39, 8)),
			21 => std_logic_vector(to_unsigned(142, 8)),
			22 => std_logic_vector(to_unsigned(199, 8)),
			23 => std_logic_vector(to_unsigned(17, 8)),
			24 => std_logic_vector(to_unsigned(187, 8)),
			25 => std_logic_vector(to_unsigned(100, 8)),
			26 => std_logic_vector(to_unsigned(1, 8)),
			27 => std_logic_vector(to_unsigned(211, 8)),
			28 => std_logic_vector(to_unsigned(118, 8)),
			29 => std_logic_vector(to_unsigned(145, 8)),
			30 => std_logic_vector(to_unsigned(37, 8)),
			31 => std_logic_vector(to_unsigned(254, 8)),
			32 => std_logic_vector(to_unsigned(187, 8)),
			33 => std_logic_vector(to_unsigned(35, 8)),
			34 => std_logic_vector(to_unsigned(63, 8)),
			35 => std_logic_vector(to_unsigned(204, 8)),
			36 => std_logic_vector(to_unsigned(215, 8)),
			37 => std_logic_vector(to_unsigned(53, 8)),
			38 => std_logic_vector(to_unsigned(62, 8)),
			39 => std_logic_vector(to_unsigned(26, 8)),
			40 => std_logic_vector(to_unsigned(101, 8)),
			41 => std_logic_vector(to_unsigned(116, 8)),
			42 => std_logic_vector(to_unsigned(42, 8)),
			43 => std_logic_vector(to_unsigned(231, 8)),
			44 => std_logic_vector(to_unsigned(46, 8)),
			45 => std_logic_vector(to_unsigned(27, 8)),
			46 => std_logic_vector(to_unsigned(137, 8)),
			47 => std_logic_vector(to_unsigned(83, 8)),
			48 => std_logic_vector(to_unsigned(20, 8)),
			49 => std_logic_vector(to_unsigned(230, 8)),
			50 => std_logic_vector(to_unsigned(51, 8)),
			51 => std_logic_vector(to_unsigned(204, 8)),
			52 => std_logic_vector(to_unsigned(228, 8)),
			53 => std_logic_vector(to_unsigned(38, 8)),
			54 => std_logic_vector(to_unsigned(112, 8)),
			55 => std_logic_vector(to_unsigned(45, 8)),
			56 => std_logic_vector(to_unsigned(139, 8)),
			57 => std_logic_vector(to_unsigned(188, 8)),
			58 => std_logic_vector(to_unsigned(168, 8)),
			59 => std_logic_vector(to_unsigned(189, 8)),
			60 => std_logic_vector(to_unsigned(109, 8)),
			61 => std_logic_vector(to_unsigned(253, 8)),
			62 => std_logic_vector(to_unsigned(234, 8)),
			63 => std_logic_vector(to_unsigned(142, 8)),
			64 => std_logic_vector(to_unsigned(67, 8)),
			65 => std_logic_vector(to_unsigned(144, 8)),
			66 => std_logic_vector(to_unsigned(56, 8)),
			67 => std_logic_vector(to_unsigned(221, 8)),
			68 => std_logic_vector(to_unsigned(40, 8)),
			69 => std_logic_vector(to_unsigned(95, 8)),
			70 => std_logic_vector(to_unsigned(80, 8)),
			71 => std_logic_vector(to_unsigned(120, 8)),
			72 => std_logic_vector(to_unsigned(80, 8)),
			73 => std_logic_vector(to_unsigned(221, 8)),
			74 => std_logic_vector(to_unsigned(69, 8)),
			75 => std_logic_vector(to_unsigned(41, 8)),
			76 => std_logic_vector(to_unsigned(21, 8)),
			77 => std_logic_vector(to_unsigned(104, 8)),
			78 => std_logic_vector(to_unsigned(123, 8)),
			79 => std_logic_vector(to_unsigned(119, 8)),
			80 => std_logic_vector(to_unsigned(221, 8)),
			81 => std_logic_vector(to_unsigned(68, 8)),
			82 => std_logic_vector(to_unsigned(106, 8)),
			83 => std_logic_vector(to_unsigned(225, 8)),
			84 => std_logic_vector(to_unsigned(103, 8)),
			85 => std_logic_vector(to_unsigned(7, 8)),
			86 => std_logic_vector(to_unsigned(188, 8)),
			87 => std_logic_vector(to_unsigned(231, 8)),
			88 => std_logic_vector(to_unsigned(121, 8)),
			89 => std_logic_vector(to_unsigned(255, 8)),
			90 => std_logic_vector(to_unsigned(140, 8)),
			91 => std_logic_vector(to_unsigned(162, 8)),
			92 => std_logic_vector(to_unsigned(30, 8)),
			93 => std_logic_vector(to_unsigned(164, 8)),
			94 => std_logic_vector(to_unsigned(195, 8)),
			95 => std_logic_vector(to_unsigned(10, 8)),
			96 => std_logic_vector(to_unsigned(132, 8)),
			97 => std_logic_vector(to_unsigned(25, 8)),
			98 => std_logic_vector(to_unsigned(254, 8)),
			99 => std_logic_vector(to_unsigned(201, 8)),
			100 => std_logic_vector(to_unsigned(211, 8)),
			101 => std_logic_vector(to_unsigned(127, 8)),
			102 => std_logic_vector(to_unsigned(138, 8)),
			103 => std_logic_vector(to_unsigned(196, 8)),
			104 => std_logic_vector(to_unsigned(114, 8)),
			105 => std_logic_vector(to_unsigned(59, 8)),
			106 => std_logic_vector(to_unsigned(160, 8)),
			107 => std_logic_vector(to_unsigned(222, 8)),
			108 => std_logic_vector(to_unsigned(205, 8)),
			109 => std_logic_vector(to_unsigned(93, 8)),
			110 => std_logic_vector(to_unsigned(38, 8)),
			111 => std_logic_vector(to_unsigned(127, 8)),
			112 => std_logic_vector(to_unsigned(169, 8)),
			113 => std_logic_vector(to_unsigned(123, 8)),
			114 => std_logic_vector(to_unsigned(230, 8)),
			115 => std_logic_vector(to_unsigned(248, 8)),
			116 => std_logic_vector(to_unsigned(194, 8)),
			117 => std_logic_vector(to_unsigned(207, 8)),
			118 => std_logic_vector(to_unsigned(47, 8)),
			119 => std_logic_vector(to_unsigned(250, 8)),
			120 => std_logic_vector(to_unsigned(205, 8)),
			121 => std_logic_vector(to_unsigned(83, 8)),
			122 => std_logic_vector(to_unsigned(255, 8)),
			123 => std_logic_vector(to_unsigned(162, 8)),
			124 => std_logic_vector(to_unsigned(143, 8)),
			125 => std_logic_vector(to_unsigned(125, 8)),
			126 => std_logic_vector(to_unsigned(45, 8)),
			127 => std_logic_vector(to_unsigned(107, 8)),
			128 => std_logic_vector(to_unsigned(105, 8)),
			129 => std_logic_vector(to_unsigned(189, 8)),
			130 => std_logic_vector(to_unsigned(199, 8)),
			131 => std_logic_vector(to_unsigned(72, 8)),
			132 => std_logic_vector(to_unsigned(124, 8)),
			133 => std_logic_vector(to_unsigned(168, 8)),
			134 => std_logic_vector(to_unsigned(11, 8)),
			135 => std_logic_vector(to_unsigned(23, 8)),
			136 => std_logic_vector(to_unsigned(61, 8)),
			137 => std_logic_vector(to_unsigned(239, 8)),
			138 => std_logic_vector(to_unsigned(177, 8)),
			139 => std_logic_vector(to_unsigned(145, 8)),
			140 => std_logic_vector(to_unsigned(112, 8)),
			141 => std_logic_vector(to_unsigned(2, 8)),
			142 => std_logic_vector(to_unsigned(52, 8)),
			143 => std_logic_vector(to_unsigned(94, 8)),
			144 => std_logic_vector(to_unsigned(83, 8)),
			145 => std_logic_vector(to_unsigned(200, 8)),
			146 => std_logic_vector(to_unsigned(0, 8)),
			147 => std_logic_vector(to_unsigned(217, 8)),
			148 => std_logic_vector(to_unsigned(183, 8)),
			149 => std_logic_vector(to_unsigned(79, 8)),
			150 => std_logic_vector(to_unsigned(34, 8)),
			151 => std_logic_vector(to_unsigned(80, 8)),
			152 => std_logic_vector(to_unsigned(7, 8)),
			153 => std_logic_vector(to_unsigned(246, 8)),
			154 => std_logic_vector(to_unsigned(118, 8)),
			155 => std_logic_vector(to_unsigned(10, 8)),
			156 => std_logic_vector(to_unsigned(238, 8)),
			157 => std_logic_vector(to_unsigned(167, 8)),
			158 => std_logic_vector(to_unsigned(28, 8)),
			159 => std_logic_vector(to_unsigned(155, 8)),
			160 => std_logic_vector(to_unsigned(74, 8)),
			161 => std_logic_vector(to_unsigned(21, 8)),
			162 => std_logic_vector(to_unsigned(182, 8)),
			163 => std_logic_vector(to_unsigned(115, 8)),
			164 => std_logic_vector(to_unsigned(52, 8)),
			165 => std_logic_vector(to_unsigned(247, 8)),
			166 => std_logic_vector(to_unsigned(245, 8)),
			167 => std_logic_vector(to_unsigned(231, 8)),
			168 => std_logic_vector(to_unsigned(107, 8)),
			169 => std_logic_vector(to_unsigned(175, 8)),
			170 => std_logic_vector(to_unsigned(70, 8)),
			171 => std_logic_vector(to_unsigned(169, 8)),
			172 => std_logic_vector(to_unsigned(115, 8)),
			173 => std_logic_vector(to_unsigned(89, 8)),
			174 => std_logic_vector(to_unsigned(16, 8)),
			175 => std_logic_vector(to_unsigned(122, 8)),
			176 => std_logic_vector(to_unsigned(132, 8)),
			177 => std_logic_vector(to_unsigned(212, 8)),
			178 => std_logic_vector(to_unsigned(142, 8)),
			179 => std_logic_vector(to_unsigned(33, 8)),
			180 => std_logic_vector(to_unsigned(25, 8)),
			181 => std_logic_vector(to_unsigned(31, 8)),
			182 => std_logic_vector(to_unsigned(225, 8)),
			183 => std_logic_vector(to_unsigned(202, 8)),
			184 => std_logic_vector(to_unsigned(8, 8)),
			185 => std_logic_vector(to_unsigned(75, 8)),
			186 => std_logic_vector(to_unsigned(103, 8)),
			187 => std_logic_vector(to_unsigned(235, 8)),
			188 => std_logic_vector(to_unsigned(0, 8)),
			189 => std_logic_vector(to_unsigned(210, 8)),
			190 => std_logic_vector(to_unsigned(29, 8)),
			191 => std_logic_vector(to_unsigned(245, 8)),
			192 => std_logic_vector(to_unsigned(71, 8)),
			193 => std_logic_vector(to_unsigned(115, 8)),
			194 => std_logic_vector(to_unsigned(235, 8)),
			195 => std_logic_vector(to_unsigned(101, 8)),
			196 => std_logic_vector(to_unsigned(93, 8)),
			197 => std_logic_vector(to_unsigned(13, 8)),
			198 => std_logic_vector(to_unsigned(27, 8)),
			199 => std_logic_vector(to_unsigned(211, 8)),
			200 => std_logic_vector(to_unsigned(25, 8)),
			201 => std_logic_vector(to_unsigned(104, 8)),
			202 => std_logic_vector(to_unsigned(145, 8)),
			203 => std_logic_vector(to_unsigned(237, 8)),
			204 => std_logic_vector(to_unsigned(190, 8)),
			205 => std_logic_vector(to_unsigned(221, 8)),
			206 => std_logic_vector(to_unsigned(12, 8)),
			207 => std_logic_vector(to_unsigned(111, 8)),
			208 => std_logic_vector(to_unsigned(18, 8)),
			209 => std_logic_vector(to_unsigned(74, 8)),
			210 => std_logic_vector(to_unsigned(113, 8)),
			211 => std_logic_vector(to_unsigned(87, 8)),
			212 => std_logic_vector(to_unsigned(74, 8)),
			213 => std_logic_vector(to_unsigned(62, 8)),
			214 => std_logic_vector(to_unsigned(149, 8)),
			215 => std_logic_vector(to_unsigned(8, 8)),
			216 => std_logic_vector(to_unsigned(94, 8)),
			217 => std_logic_vector(to_unsigned(200, 8)),
			218 => std_logic_vector(to_unsigned(157, 8)),
			219 => std_logic_vector(to_unsigned(157, 8)),
			220 => std_logic_vector(to_unsigned(40, 8)),
			221 => std_logic_vector(to_unsigned(79, 8)),
			222 => std_logic_vector(to_unsigned(163, 8)),
			223 => std_logic_vector(to_unsigned(131, 8)),
			224 => std_logic_vector(to_unsigned(60, 8)),
			225 => std_logic_vector(to_unsigned(8, 8)),
			226 => std_logic_vector(to_unsigned(244, 8)),
			227 => std_logic_vector(to_unsigned(142, 8)),
			228 => std_logic_vector(to_unsigned(143, 8)),
			229 => std_logic_vector(to_unsigned(195, 8)),
			230 => std_logic_vector(to_unsigned(0, 8)),
			231 => std_logic_vector(to_unsigned(202, 8)),
			232 => std_logic_vector(to_unsigned(232, 8)),
			233 => std_logic_vector(to_unsigned(176, 8)),
			234 => std_logic_vector(to_unsigned(7, 8)),
			235 => std_logic_vector(to_unsigned(156, 8)),
			236 => std_logic_vector(to_unsigned(244, 8)),
			237 => std_logic_vector(to_unsigned(192, 8)),
			238 => std_logic_vector(to_unsigned(148, 8)),
			239 => std_logic_vector(to_unsigned(93, 8)),
			240 => std_logic_vector(to_unsigned(100, 8)),
			241 => std_logic_vector(to_unsigned(95, 8)),
			242 => std_logic_vector(to_unsigned(192, 8)),
			243 => std_logic_vector(to_unsigned(99, 8)),
			244 => std_logic_vector(to_unsigned(27, 8)),
			245 => std_logic_vector(to_unsigned(166, 8)),
			246 => std_logic_vector(to_unsigned(45, 8)),
			247 => std_logic_vector(to_unsigned(82, 8)),
			248 => std_logic_vector(to_unsigned(95, 8)),
			249 => std_logic_vector(to_unsigned(166, 8)),
			250 => std_logic_vector(to_unsigned(122, 8)),
			251 => std_logic_vector(to_unsigned(100, 8)),
			252 => std_logic_vector(to_unsigned(154, 8)),
			253 => std_logic_vector(to_unsigned(163, 8)),
			254 => std_logic_vector(to_unsigned(107, 8)),
			255 => std_logic_vector(to_unsigned(147, 8)),
			256 => std_logic_vector(to_unsigned(59, 8)),
			257 => std_logic_vector(to_unsigned(4, 8)),
			258 => std_logic_vector(to_unsigned(165, 8)),
			259 => std_logic_vector(to_unsigned(149, 8)),
			260 => std_logic_vector(to_unsigned(9, 8)),
			261 => std_logic_vector(to_unsigned(11, 8)),
			262 => std_logic_vector(to_unsigned(137, 8)),
			263 => std_logic_vector(to_unsigned(198, 8)),
			264 => std_logic_vector(to_unsigned(244, 8)),
			265 => std_logic_vector(to_unsigned(166, 8)),
			266 => std_logic_vector(to_unsigned(203, 8)),
			267 => std_logic_vector(to_unsigned(196, 8)),
			268 => std_logic_vector(to_unsigned(184, 8)),
			269 => std_logic_vector(to_unsigned(63, 8)),
			270 => std_logic_vector(to_unsigned(30, 8)),
			271 => std_logic_vector(to_unsigned(133, 8)),
			272 => std_logic_vector(to_unsigned(97, 8)),
			273 => std_logic_vector(to_unsigned(25, 8)),
			274 => std_logic_vector(to_unsigned(230, 8)),
			275 => std_logic_vector(to_unsigned(179, 8)),
			276 => std_logic_vector(to_unsigned(63, 8)),
			277 => std_logic_vector(to_unsigned(255, 8)),
			278 => std_logic_vector(to_unsigned(1, 8)),
			279 => std_logic_vector(to_unsigned(210, 8)),
			280 => std_logic_vector(to_unsigned(26, 8)),
			281 => std_logic_vector(to_unsigned(202, 8)),
			282 => std_logic_vector(to_unsigned(52, 8)),
			283 => std_logic_vector(to_unsigned(5, 8)),
			284 => std_logic_vector(to_unsigned(40, 8)),
			285 => std_logic_vector(to_unsigned(107, 8)),
			286 => std_logic_vector(to_unsigned(213, 8)),
			287 => std_logic_vector(to_unsigned(66, 8)),
			288 => std_logic_vector(to_unsigned(156, 8)),
			289 => std_logic_vector(to_unsigned(210, 8)),
			290 => std_logic_vector(to_unsigned(23, 8)),
			291 => std_logic_vector(to_unsigned(130, 8)),
			292 => std_logic_vector(to_unsigned(4, 8)),
			293 => std_logic_vector(to_unsigned(207, 8)),
			294 => std_logic_vector(to_unsigned(144, 8)),
			295 => std_logic_vector(to_unsigned(232, 8)),
			296 => std_logic_vector(to_unsigned(37, 8)),
			297 => std_logic_vector(to_unsigned(106, 8)),
			298 => std_logic_vector(to_unsigned(45, 8)),
			299 => std_logic_vector(to_unsigned(106, 8)),
			300 => std_logic_vector(to_unsigned(24, 8)),
			301 => std_logic_vector(to_unsigned(26, 8)),
			302 => std_logic_vector(to_unsigned(163, 8)),
			303 => std_logic_vector(to_unsigned(219, 8)),
			304 => std_logic_vector(to_unsigned(211, 8)),
			305 => std_logic_vector(to_unsigned(39, 8)),
			306 => std_logic_vector(to_unsigned(39, 8)),
			307 => std_logic_vector(to_unsigned(135, 8)),
			308 => std_logic_vector(to_unsigned(217, 8)),
			309 => std_logic_vector(to_unsigned(106, 8)),
			310 => std_logic_vector(to_unsigned(17, 8)),
			311 => std_logic_vector(to_unsigned(247, 8)),
			312 => std_logic_vector(to_unsigned(188, 8)),
			313 => std_logic_vector(to_unsigned(98, 8)),
			314 => std_logic_vector(to_unsigned(119, 8)),
			315 => std_logic_vector(to_unsigned(68, 8)),
			316 => std_logic_vector(to_unsigned(128, 8)),
			317 => std_logic_vector(to_unsigned(164, 8)),
			318 => std_logic_vector(to_unsigned(49, 8)),
			319 => std_logic_vector(to_unsigned(13, 8)),
			320 => std_logic_vector(to_unsigned(40, 8)),
			321 => std_logic_vector(to_unsigned(208, 8)),
			322 => std_logic_vector(to_unsigned(49, 8)),
			323 => std_logic_vector(to_unsigned(45, 8)),
			324 => std_logic_vector(to_unsigned(15, 8)),
			325 => std_logic_vector(to_unsigned(154, 8)),
			326 => std_logic_vector(to_unsigned(218, 8)),
			327 => std_logic_vector(to_unsigned(103, 8)),
			328 => std_logic_vector(to_unsigned(254, 8)),
			329 => std_logic_vector(to_unsigned(124, 8)),
			330 => std_logic_vector(to_unsigned(182, 8)),
			331 => std_logic_vector(to_unsigned(15, 8)),
			332 => std_logic_vector(to_unsigned(233, 8)),
			333 => std_logic_vector(to_unsigned(165, 8)),
			334 => std_logic_vector(to_unsigned(114, 8)),
			335 => std_logic_vector(to_unsigned(115, 8)),
			336 => std_logic_vector(to_unsigned(220, 8)),
			337 => std_logic_vector(to_unsigned(96, 8)),
			338 => std_logic_vector(to_unsigned(247, 8)),
			339 => std_logic_vector(to_unsigned(187, 8)),
			340 => std_logic_vector(to_unsigned(133, 8)),
			341 => std_logic_vector(to_unsigned(95, 8)),
			342 => std_logic_vector(to_unsigned(237, 8)),
			343 => std_logic_vector(to_unsigned(109, 8)),
			344 => std_logic_vector(to_unsigned(229, 8)),
			345 => std_logic_vector(to_unsigned(43, 8)),
			346 => std_logic_vector(to_unsigned(190, 8)),
			347 => std_logic_vector(to_unsigned(185, 8)),
			348 => std_logic_vector(to_unsigned(123, 8)),
			349 => std_logic_vector(to_unsigned(46, 8)),
			350 => std_logic_vector(to_unsigned(78, 8)),
			351 => std_logic_vector(to_unsigned(18, 8)),
			352 => std_logic_vector(to_unsigned(90, 8)),
			353 => std_logic_vector(to_unsigned(150, 8)),
			354 => std_logic_vector(to_unsigned(98, 8)),
			355 => std_logic_vector(to_unsigned(50, 8)),
			356 => std_logic_vector(to_unsigned(201, 8)),
			357 => std_logic_vector(to_unsigned(13, 8)),
			358 => std_logic_vector(to_unsigned(66, 8)),
			359 => std_logic_vector(to_unsigned(81, 8)),
			360 => std_logic_vector(to_unsigned(70, 8)),
			361 => std_logic_vector(to_unsigned(32, 8)),
			362 => std_logic_vector(to_unsigned(37, 8)),
			363 => std_logic_vector(to_unsigned(243, 8)),
			364 => std_logic_vector(to_unsigned(180, 8)),
			365 => std_logic_vector(to_unsigned(17, 8)),
			366 => std_logic_vector(to_unsigned(138, 8)),
			367 => std_logic_vector(to_unsigned(7, 8)),
			368 => std_logic_vector(to_unsigned(248, 8)),
			369 => std_logic_vector(to_unsigned(96, 8)),
			370 => std_logic_vector(to_unsigned(201, 8)),
			371 => std_logic_vector(to_unsigned(194, 8)),
			372 => std_logic_vector(to_unsigned(252, 8)),
			373 => std_logic_vector(to_unsigned(154, 8)),
			374 => std_logic_vector(to_unsigned(109, 8)),
			375 => std_logic_vector(to_unsigned(149, 8)),
			376 => std_logic_vector(to_unsigned(243, 8)),
			377 => std_logic_vector(to_unsigned(32, 8)),
			378 => std_logic_vector(to_unsigned(187, 8)),
			379 => std_logic_vector(to_unsigned(195, 8)),
			380 => std_logic_vector(to_unsigned(15, 8)),
			381 => std_logic_vector(to_unsigned(97, 8)),
			382 => std_logic_vector(to_unsigned(162, 8)),
			383 => std_logic_vector(to_unsigned(207, 8)),
			384 => std_logic_vector(to_unsigned(8, 8)),
			385 => std_logic_vector(to_unsigned(238, 8)),
			386 => std_logic_vector(to_unsigned(175, 8)),
			387 => std_logic_vector(to_unsigned(104, 8)),
			388 => std_logic_vector(to_unsigned(124, 8)),
			389 => std_logic_vector(to_unsigned(127, 8)),
			390 => std_logic_vector(to_unsigned(225, 8)),
			391 => std_logic_vector(to_unsigned(25, 8)),
			392 => std_logic_vector(to_unsigned(198, 8)),
			393 => std_logic_vector(to_unsigned(197, 8)),
			394 => std_logic_vector(to_unsigned(14, 8)),
			395 => std_logic_vector(to_unsigned(45, 8)),
			396 => std_logic_vector(to_unsigned(121, 8)),
			397 => std_logic_vector(to_unsigned(246, 8)),
			398 => std_logic_vector(to_unsigned(222, 8)),
			399 => std_logic_vector(to_unsigned(186, 8)),
			400 => std_logic_vector(to_unsigned(165, 8)),
			401 => std_logic_vector(to_unsigned(12, 8)),
			402 => std_logic_vector(to_unsigned(170, 8)),
			403 => std_logic_vector(to_unsigned(24, 8)),
			404 => std_logic_vector(to_unsigned(4, 8)),
			405 => std_logic_vector(to_unsigned(11, 8)),
			406 => std_logic_vector(to_unsigned(20, 8)),
			407 => std_logic_vector(to_unsigned(50, 8)),
			408 => std_logic_vector(to_unsigned(27, 8)),
			409 => std_logic_vector(to_unsigned(158, 8)),
			410 => std_logic_vector(to_unsigned(92, 8)),
			411 => std_logic_vector(to_unsigned(191, 8)),
			412 => std_logic_vector(to_unsigned(210, 8)),
			413 => std_logic_vector(to_unsigned(21, 8)),
			414 => std_logic_vector(to_unsigned(188, 8)),
			415 => std_logic_vector(to_unsigned(36, 8)),
			416 => std_logic_vector(to_unsigned(56, 8)),
			417 => std_logic_vector(to_unsigned(86, 8)),
			418 => std_logic_vector(to_unsigned(52, 8)),
			419 => std_logic_vector(to_unsigned(106, 8)),
			420 => std_logic_vector(to_unsigned(120, 8)),
			421 => std_logic_vector(to_unsigned(236, 8)),
			422 => std_logic_vector(to_unsigned(202, 8)),
			423 => std_logic_vector(to_unsigned(92, 8)),
			424 => std_logic_vector(to_unsigned(172, 8)),
			425 => std_logic_vector(to_unsigned(196, 8)),
			426 => std_logic_vector(to_unsigned(242, 8)),
			427 => std_logic_vector(to_unsigned(41, 8)),
			428 => std_logic_vector(to_unsigned(255, 8)),
			429 => std_logic_vector(to_unsigned(255, 8)),
			430 => std_logic_vector(to_unsigned(197, 8)),
			431 => std_logic_vector(to_unsigned(3, 8)),
			432 => std_logic_vector(to_unsigned(241, 8)),
			433 => std_logic_vector(to_unsigned(234, 8)),
			434 => std_logic_vector(to_unsigned(20, 8)),
			435 => std_logic_vector(to_unsigned(156, 8)),
			436 => std_logic_vector(to_unsigned(186, 8)),
			437 => std_logic_vector(to_unsigned(142, 8)),
			438 => std_logic_vector(to_unsigned(80, 8)),
			439 => std_logic_vector(to_unsigned(28, 8)),
			440 => std_logic_vector(to_unsigned(45, 8)),
			441 => std_logic_vector(to_unsigned(103, 8)),
			442 => std_logic_vector(to_unsigned(58, 8)),
			443 => std_logic_vector(to_unsigned(27, 8)),
			444 => std_logic_vector(to_unsigned(66, 8)),
			445 => std_logic_vector(to_unsigned(54, 8)),
			446 => std_logic_vector(to_unsigned(40, 8)),
			447 => std_logic_vector(to_unsigned(49, 8)),
			448 => std_logic_vector(to_unsigned(147, 8)),
			449 => std_logic_vector(to_unsigned(184, 8)),
			450 => std_logic_vector(to_unsigned(100, 8)),
			451 => std_logic_vector(to_unsigned(53, 8)),
			452 => std_logic_vector(to_unsigned(126, 8)),
			453 => std_logic_vector(to_unsigned(26, 8)),
			454 => std_logic_vector(to_unsigned(53, 8)),
			455 => std_logic_vector(to_unsigned(90, 8)),
			456 => std_logic_vector(to_unsigned(16, 8)),
			457 => std_logic_vector(to_unsigned(225, 8)),
			458 => std_logic_vector(to_unsigned(191, 8)),
			459 => std_logic_vector(to_unsigned(182, 8)),
			460 => std_logic_vector(to_unsigned(86, 8)),
			461 => std_logic_vector(to_unsigned(102, 8)),
			462 => std_logic_vector(to_unsigned(234, 8)),
			463 => std_logic_vector(to_unsigned(138, 8)),
			464 => std_logic_vector(to_unsigned(250, 8)),
			465 => std_logic_vector(to_unsigned(210, 8)),
			466 => std_logic_vector(to_unsigned(128, 8)),
			467 => std_logic_vector(to_unsigned(0, 8)),
			468 => std_logic_vector(to_unsigned(160, 8)),
			469 => std_logic_vector(to_unsigned(200, 8)),
			470 => std_logic_vector(to_unsigned(198, 8)),
			471 => std_logic_vector(to_unsigned(63, 8)),
			472 => std_logic_vector(to_unsigned(40, 8)),
			473 => std_logic_vector(to_unsigned(216, 8)),
			474 => std_logic_vector(to_unsigned(52, 8)),
			475 => std_logic_vector(to_unsigned(62, 8)),
			476 => std_logic_vector(to_unsigned(205, 8)),
			477 => std_logic_vector(to_unsigned(75, 8)),
			478 => std_logic_vector(to_unsigned(41, 8)),
			479 => std_logic_vector(to_unsigned(128, 8)),
			480 => std_logic_vector(to_unsigned(64, 8)),
			481 => std_logic_vector(to_unsigned(204, 8)),
			482 => std_logic_vector(to_unsigned(194, 8)),
			483 => std_logic_vector(to_unsigned(255, 8)),
			484 => std_logic_vector(to_unsigned(63, 8)),
			485 => std_logic_vector(to_unsigned(134, 8)),
			486 => std_logic_vector(to_unsigned(7, 8)),
			487 => std_logic_vector(to_unsigned(159, 8)),
			488 => std_logic_vector(to_unsigned(161, 8)),
			489 => std_logic_vector(to_unsigned(107, 8)),
			490 => std_logic_vector(to_unsigned(237, 8)),
			491 => std_logic_vector(to_unsigned(47, 8)),
			492 => std_logic_vector(to_unsigned(106, 8)),
			493 => std_logic_vector(to_unsigned(158, 8)),
			494 => std_logic_vector(to_unsigned(132, 8)),
			495 => std_logic_vector(to_unsigned(55, 8)),
			496 => std_logic_vector(to_unsigned(123, 8)),
			497 => std_logic_vector(to_unsigned(158, 8)),
			498 => std_logic_vector(to_unsigned(138, 8)),
			499 => std_logic_vector(to_unsigned(170, 8)),
			500 => std_logic_vector(to_unsigned(237, 8)),
			501 => std_logic_vector(to_unsigned(113, 8)),
			502 => std_logic_vector(to_unsigned(68, 8)),
			503 => std_logic_vector(to_unsigned(111, 8)),
			504 => std_logic_vector(to_unsigned(230, 8)),
			505 => std_logic_vector(to_unsigned(63, 8)),
			506 => std_logic_vector(to_unsigned(244, 8)),
			507 => std_logic_vector(to_unsigned(181, 8)),
			508 => std_logic_vector(to_unsigned(213, 8)),
			509 => std_logic_vector(to_unsigned(39, 8)),
			510 => std_logic_vector(to_unsigned(199, 8)),
			511 => std_logic_vector(to_unsigned(141, 8)),
			512 => std_logic_vector(to_unsigned(76, 8)),
			513 => std_logic_vector(to_unsigned(226, 8)),
			514 => std_logic_vector(to_unsigned(64, 8)),
			515 => std_logic_vector(to_unsigned(123, 8)),
			516 => std_logic_vector(to_unsigned(17, 8)),
			517 => std_logic_vector(to_unsigned(136, 8)),
			518 => std_logic_vector(to_unsigned(134, 8)),
			519 => std_logic_vector(to_unsigned(241, 8)),
			520 => std_logic_vector(to_unsigned(112, 8)),
			521 => std_logic_vector(to_unsigned(152, 8)),
			522 => std_logic_vector(to_unsigned(72, 8)),
			523 => std_logic_vector(to_unsigned(95, 8)),
			524 => std_logic_vector(to_unsigned(173, 8)),
			525 => std_logic_vector(to_unsigned(83, 8)),
			526 => std_logic_vector(to_unsigned(2, 8)),
			527 => std_logic_vector(to_unsigned(106, 8)),
			528 => std_logic_vector(to_unsigned(69, 8)),
			529 => std_logic_vector(to_unsigned(63, 8)),
			530 => std_logic_vector(to_unsigned(74, 8)),
			531 => std_logic_vector(to_unsigned(99, 8)),
			532 => std_logic_vector(to_unsigned(227, 8)),
			533 => std_logic_vector(to_unsigned(101, 8)),
			534 => std_logic_vector(to_unsigned(209, 8)),
			535 => std_logic_vector(to_unsigned(158, 8)),
			536 => std_logic_vector(to_unsigned(62, 8)),
			537 => std_logic_vector(to_unsigned(147, 8)),
			538 => std_logic_vector(to_unsigned(32, 8)),
			539 => std_logic_vector(to_unsigned(134, 8)),
			540 => std_logic_vector(to_unsigned(116, 8)),
			541 => std_logic_vector(to_unsigned(150, 8)),
			542 => std_logic_vector(to_unsigned(187, 8)),
			543 => std_logic_vector(to_unsigned(128, 8)),
			544 => std_logic_vector(to_unsigned(117, 8)),
			545 => std_logic_vector(to_unsigned(5, 8)),
			546 => std_logic_vector(to_unsigned(143, 8)),
			547 => std_logic_vector(to_unsigned(229, 8)),
			548 => std_logic_vector(to_unsigned(118, 8)),
			549 => std_logic_vector(to_unsigned(144, 8)),
			550 => std_logic_vector(to_unsigned(184, 8)),
			551 => std_logic_vector(to_unsigned(112, 8)),
			552 => std_logic_vector(to_unsigned(156, 8)),
			553 => std_logic_vector(to_unsigned(65, 8)),
			554 => std_logic_vector(to_unsigned(8, 8)),
			555 => std_logic_vector(to_unsigned(62, 8)),
			556 => std_logic_vector(to_unsigned(73, 8)),
			557 => std_logic_vector(to_unsigned(197, 8)),
			558 => std_logic_vector(to_unsigned(90, 8)),
			559 => std_logic_vector(to_unsigned(167, 8)),
			560 => std_logic_vector(to_unsigned(66, 8)),
			561 => std_logic_vector(to_unsigned(97, 8)),
			562 => std_logic_vector(to_unsigned(130, 8)),
			563 => std_logic_vector(to_unsigned(108, 8)),
			564 => std_logic_vector(to_unsigned(184, 8)),
			565 => std_logic_vector(to_unsigned(190, 8)),
			566 => std_logic_vector(to_unsigned(226, 8)),
			567 => std_logic_vector(to_unsigned(61, 8)),
			568 => std_logic_vector(to_unsigned(24, 8)),
			569 => std_logic_vector(to_unsigned(124, 8)),
			570 => std_logic_vector(to_unsigned(164, 8)),
			571 => std_logic_vector(to_unsigned(241, 8)),
			572 => std_logic_vector(to_unsigned(50, 8)),
			573 => std_logic_vector(to_unsigned(69, 8)),
			574 => std_logic_vector(to_unsigned(57, 8)),
			575 => std_logic_vector(to_unsigned(129, 8)),
			576 => std_logic_vector(to_unsigned(43, 8)),
			577 => std_logic_vector(to_unsigned(175, 8)),
			578 => std_logic_vector(to_unsigned(179, 8)),
			579 => std_logic_vector(to_unsigned(214, 8)),
			580 => std_logic_vector(to_unsigned(203, 8)),
			581 => std_logic_vector(to_unsigned(37, 8)),
			582 => std_logic_vector(to_unsigned(244, 8)),
			583 => std_logic_vector(to_unsigned(232, 8)),
			584 => std_logic_vector(to_unsigned(120, 8)),
			585 => std_logic_vector(to_unsigned(114, 8)),
			586 => std_logic_vector(to_unsigned(15, 8)),
			587 => std_logic_vector(to_unsigned(187, 8)),
			588 => std_logic_vector(to_unsigned(115, 8)),
			589 => std_logic_vector(to_unsigned(51, 8)),
			590 => std_logic_vector(to_unsigned(1, 8)),
			591 => std_logic_vector(to_unsigned(75, 8)),
			592 => std_logic_vector(to_unsigned(95, 8)),
			593 => std_logic_vector(to_unsigned(113, 8)),
			594 => std_logic_vector(to_unsigned(242, 8)),
			595 => std_logic_vector(to_unsigned(36, 8)),
			596 => std_logic_vector(to_unsigned(86, 8)),
			597 => std_logic_vector(to_unsigned(37, 8)),
			598 => std_logic_vector(to_unsigned(118, 8)),
			599 => std_logic_vector(to_unsigned(17, 8)),
			600 => std_logic_vector(to_unsigned(253, 8)),
			601 => std_logic_vector(to_unsigned(173, 8)),
			602 => std_logic_vector(to_unsigned(146, 8)),
			603 => std_logic_vector(to_unsigned(83, 8)),
			604 => std_logic_vector(to_unsigned(84, 8)),
			605 => std_logic_vector(to_unsigned(79, 8)),
			606 => std_logic_vector(to_unsigned(83, 8)),
			607 => std_logic_vector(to_unsigned(55, 8)),
			608 => std_logic_vector(to_unsigned(99, 8)),
			609 => std_logic_vector(to_unsigned(139, 8)),
			610 => std_logic_vector(to_unsigned(214, 8)),
			611 => std_logic_vector(to_unsigned(84, 8)),
			612 => std_logic_vector(to_unsigned(172, 8)),
			613 => std_logic_vector(to_unsigned(162, 8)),
			614 => std_logic_vector(to_unsigned(66, 8)),
			615 => std_logic_vector(to_unsigned(137, 8)),
			616 => std_logic_vector(to_unsigned(188, 8)),
			617 => std_logic_vector(to_unsigned(80, 8)),
			618 => std_logic_vector(to_unsigned(132, 8)),
			619 => std_logic_vector(to_unsigned(33, 8)),
			620 => std_logic_vector(to_unsigned(195, 8)),
			621 => std_logic_vector(to_unsigned(73, 8)),
			622 => std_logic_vector(to_unsigned(194, 8)),
			623 => std_logic_vector(to_unsigned(25, 8)),
			624 => std_logic_vector(to_unsigned(36, 8)),
			625 => std_logic_vector(to_unsigned(44, 8)),
			626 => std_logic_vector(to_unsigned(183, 8)),
			627 => std_logic_vector(to_unsigned(24, 8)),
			628 => std_logic_vector(to_unsigned(59, 8)),
			629 => std_logic_vector(to_unsigned(242, 8)),
			630 => std_logic_vector(to_unsigned(57, 8)),
			631 => std_logic_vector(to_unsigned(20, 8)),
			632 => std_logic_vector(to_unsigned(107, 8)),
			633 => std_logic_vector(to_unsigned(61, 8)),
			634 => std_logic_vector(to_unsigned(122, 8)),
			635 => std_logic_vector(to_unsigned(69, 8)),
			636 => std_logic_vector(to_unsigned(137, 8)),
			637 => std_logic_vector(to_unsigned(117, 8)),
			638 => std_logic_vector(to_unsigned(241, 8)),
			639 => std_logic_vector(to_unsigned(212, 8)),
			640 => std_logic_vector(to_unsigned(64, 8)),
			641 => std_logic_vector(to_unsigned(71, 8)),
			642 => std_logic_vector(to_unsigned(11, 8)),
			643 => std_logic_vector(to_unsigned(40, 8)),
			644 => std_logic_vector(to_unsigned(39, 8)),
			645 => std_logic_vector(to_unsigned(228, 8)),
			646 => std_logic_vector(to_unsigned(109, 8)),
			647 => std_logic_vector(to_unsigned(164, 8)),
			648 => std_logic_vector(to_unsigned(121, 8)),
			649 => std_logic_vector(to_unsigned(10, 8)),
			650 => std_logic_vector(to_unsigned(73, 8)),
			651 => std_logic_vector(to_unsigned(60, 8)),
			652 => std_logic_vector(to_unsigned(128, 8)),
			653 => std_logic_vector(to_unsigned(179, 8)),
			654 => std_logic_vector(to_unsigned(98, 8)),
			655 => std_logic_vector(to_unsigned(212, 8)),
			656 => std_logic_vector(to_unsigned(201, 8)),
			657 => std_logic_vector(to_unsigned(191, 8)),
			658 => std_logic_vector(to_unsigned(52, 8)),
			659 => std_logic_vector(to_unsigned(8, 8)),
			660 => std_logic_vector(to_unsigned(146, 8)),
			661 => std_logic_vector(to_unsigned(135, 8)),
			662 => std_logic_vector(to_unsigned(3, 8)),
			663 => std_logic_vector(to_unsigned(19, 8)),
			664 => std_logic_vector(to_unsigned(136, 8)),
			665 => std_logic_vector(to_unsigned(28, 8)),
			666 => std_logic_vector(to_unsigned(18, 8)),
			667 => std_logic_vector(to_unsigned(93, 8)),
			668 => std_logic_vector(to_unsigned(213, 8)),
			669 => std_logic_vector(to_unsigned(143, 8)),
			670 => std_logic_vector(to_unsigned(166, 8)),
			671 => std_logic_vector(to_unsigned(139, 8)),
			672 => std_logic_vector(to_unsigned(131, 8)),
			673 => std_logic_vector(to_unsigned(248, 8)),
			674 => std_logic_vector(to_unsigned(172, 8)),
			675 => std_logic_vector(to_unsigned(35, 8)),
			676 => std_logic_vector(to_unsigned(244, 8)),
			677 => std_logic_vector(to_unsigned(68, 8)),
			678 => std_logic_vector(to_unsigned(64, 8)),
			679 => std_logic_vector(to_unsigned(17, 8)),
			680 => std_logic_vector(to_unsigned(132, 8)),
			681 => std_logic_vector(to_unsigned(177, 8)),
			682 => std_logic_vector(to_unsigned(204, 8)),
			683 => std_logic_vector(to_unsigned(87, 8)),
			684 => std_logic_vector(to_unsigned(122, 8)),
			685 => std_logic_vector(to_unsigned(14, 8)),
			686 => std_logic_vector(to_unsigned(235, 8)),
			687 => std_logic_vector(to_unsigned(243, 8)),
			688 => std_logic_vector(to_unsigned(3, 8)),
			689 => std_logic_vector(to_unsigned(69, 8)),
			690 => std_logic_vector(to_unsigned(24, 8)),
			691 => std_logic_vector(to_unsigned(231, 8)),
			692 => std_logic_vector(to_unsigned(108, 8)),
			693 => std_logic_vector(to_unsigned(177, 8)),
			694 => std_logic_vector(to_unsigned(255, 8)),
			695 => std_logic_vector(to_unsigned(111, 8)),
			696 => std_logic_vector(to_unsigned(198, 8)),
			697 => std_logic_vector(to_unsigned(185, 8)),
			698 => std_logic_vector(to_unsigned(149, 8)),
			699 => std_logic_vector(to_unsigned(189, 8)),
			700 => std_logic_vector(to_unsigned(33, 8)),
			701 => std_logic_vector(to_unsigned(214, 8)),
			702 => std_logic_vector(to_unsigned(162, 8)),
			703 => std_logic_vector(to_unsigned(26, 8)),
			704 => std_logic_vector(to_unsigned(203, 8)),
			705 => std_logic_vector(to_unsigned(210, 8)),
			706 => std_logic_vector(to_unsigned(55, 8)),
			707 => std_logic_vector(to_unsigned(252, 8)),
			708 => std_logic_vector(to_unsigned(222, 8)),
			709 => std_logic_vector(to_unsigned(115, 8)),
			710 => std_logic_vector(to_unsigned(142, 8)),
			711 => std_logic_vector(to_unsigned(69, 8)),
			712 => std_logic_vector(to_unsigned(8, 8)),
			713 => std_logic_vector(to_unsigned(87, 8)),
			714 => std_logic_vector(to_unsigned(188, 8)),
			715 => std_logic_vector(to_unsigned(34, 8)),
			716 => std_logic_vector(to_unsigned(149, 8)),
			717 => std_logic_vector(to_unsigned(95, 8)),
			718 => std_logic_vector(to_unsigned(103, 8)),
			719 => std_logic_vector(to_unsigned(231, 8)),
			720 => std_logic_vector(to_unsigned(99, 8)),
			721 => std_logic_vector(to_unsigned(4, 8)),
			722 => std_logic_vector(to_unsigned(216, 8)),
			723 => std_logic_vector(to_unsigned(63, 8)),
			724 => std_logic_vector(to_unsigned(160, 8)),
			725 => std_logic_vector(to_unsigned(205, 8)),
			726 => std_logic_vector(to_unsigned(200, 8)),
			727 => std_logic_vector(to_unsigned(182, 8)),
			728 => std_logic_vector(to_unsigned(249, 8)),
			729 => std_logic_vector(to_unsigned(59, 8)),
			730 => std_logic_vector(to_unsigned(172, 8)),
			731 => std_logic_vector(to_unsigned(82, 8)),
			732 => std_logic_vector(to_unsigned(245, 8)),
			733 => std_logic_vector(to_unsigned(73, 8)),
			734 => std_logic_vector(to_unsigned(230, 8)),
			735 => std_logic_vector(to_unsigned(233, 8)),
			736 => std_logic_vector(to_unsigned(132, 8)),
			737 => std_logic_vector(to_unsigned(170, 8)),
			738 => std_logic_vector(to_unsigned(22, 8)),
			739 => std_logic_vector(to_unsigned(29, 8)),
			740 => std_logic_vector(to_unsigned(86, 8)),
			741 => std_logic_vector(to_unsigned(104, 8)),
			742 => std_logic_vector(to_unsigned(125, 8)),
			743 => std_logic_vector(to_unsigned(206, 8)),
			744 => std_logic_vector(to_unsigned(191, 8)),
			745 => std_logic_vector(to_unsigned(239, 8)),
			746 => std_logic_vector(to_unsigned(219, 8)),
			747 => std_logic_vector(to_unsigned(53, 8)),
			748 => std_logic_vector(to_unsigned(166, 8)),
			749 => std_logic_vector(to_unsigned(197, 8)),
			750 => std_logic_vector(to_unsigned(68, 8)),
			751 => std_logic_vector(to_unsigned(35, 8)),
			752 => std_logic_vector(to_unsigned(19, 8)),
			753 => std_logic_vector(to_unsigned(255, 8)),
			754 => std_logic_vector(to_unsigned(246, 8)),
			755 => std_logic_vector(to_unsigned(80, 8)),
			756 => std_logic_vector(to_unsigned(148, 8)),
			757 => std_logic_vector(to_unsigned(151, 8)),
			758 => std_logic_vector(to_unsigned(197, 8)),
			759 => std_logic_vector(to_unsigned(72, 8)),
			760 => std_logic_vector(to_unsigned(174, 8)),
			761 => std_logic_vector(to_unsigned(206, 8)),
			762 => std_logic_vector(to_unsigned(149, 8)),
			763 => std_logic_vector(to_unsigned(95, 8)),
			764 => std_logic_vector(to_unsigned(8, 8)),
			765 => std_logic_vector(to_unsigned(147, 8)),
			766 => std_logic_vector(to_unsigned(61, 8)),
			767 => std_logic_vector(to_unsigned(167, 8)),
			768 => std_logic_vector(to_unsigned(52, 8)),
			769 => std_logic_vector(to_unsigned(205, 8)),
			770 => std_logic_vector(to_unsigned(207, 8)),
			771 => std_logic_vector(to_unsigned(84, 8)),
			772 => std_logic_vector(to_unsigned(251, 8)),
			773 => std_logic_vector(to_unsigned(144, 8)),
			774 => std_logic_vector(to_unsigned(13, 8)),
			775 => std_logic_vector(to_unsigned(184, 8)),
			776 => std_logic_vector(to_unsigned(11, 8)),
			777 => std_logic_vector(to_unsigned(196, 8)),
			778 => std_logic_vector(to_unsigned(19, 8)),
			779 => std_logic_vector(to_unsigned(145, 8)),
			780 => std_logic_vector(to_unsigned(179, 8)),
			781 => std_logic_vector(to_unsigned(23, 8)),
			782 => std_logic_vector(to_unsigned(143, 8)),
			783 => std_logic_vector(to_unsigned(221, 8)),
			784 => std_logic_vector(to_unsigned(104, 8)),
			785 => std_logic_vector(to_unsigned(58, 8)),
			786 => std_logic_vector(to_unsigned(161, 8)),
			787 => std_logic_vector(to_unsigned(235, 8)),
			788 => std_logic_vector(to_unsigned(27, 8)),
			789 => std_logic_vector(to_unsigned(131, 8)),
			790 => std_logic_vector(to_unsigned(85, 8)),
			791 => std_logic_vector(to_unsigned(34, 8)),
			792 => std_logic_vector(to_unsigned(123, 8)),
			793 => std_logic_vector(to_unsigned(251, 8)),
			794 => std_logic_vector(to_unsigned(66, 8)),
			795 => std_logic_vector(to_unsigned(167, 8)),
			796 => std_logic_vector(to_unsigned(77, 8)),
			797 => std_logic_vector(to_unsigned(83, 8)),
			798 => std_logic_vector(to_unsigned(216, 8)),
			799 => std_logic_vector(to_unsigned(89, 8)),
			800 => std_logic_vector(to_unsigned(209, 8)),
			801 => std_logic_vector(to_unsigned(122, 8)),
			802 => std_logic_vector(to_unsigned(183, 8)),
			803 => std_logic_vector(to_unsigned(115, 8)),
			804 => std_logic_vector(to_unsigned(0, 8)),
			805 => std_logic_vector(to_unsigned(183, 8)),
			806 => std_logic_vector(to_unsigned(48, 8)),
			807 => std_logic_vector(to_unsigned(254, 8)),
			808 => std_logic_vector(to_unsigned(20, 8)),
			809 => std_logic_vector(to_unsigned(84, 8)),
			810 => std_logic_vector(to_unsigned(191, 8)),
			811 => std_logic_vector(to_unsigned(94, 8)),
			812 => std_logic_vector(to_unsigned(62, 8)),
			813 => std_logic_vector(to_unsigned(199, 8)),
			814 => std_logic_vector(to_unsigned(156, 8)),
			815 => std_logic_vector(to_unsigned(72, 8)),
			816 => std_logic_vector(to_unsigned(242, 8)),
			817 => std_logic_vector(to_unsigned(181, 8)),
			818 => std_logic_vector(to_unsigned(87, 8)),
			819 => std_logic_vector(to_unsigned(26, 8)),
			820 => std_logic_vector(to_unsigned(121, 8)),
			821 => std_logic_vector(to_unsigned(25, 8)),
			822 => std_logic_vector(to_unsigned(60, 8)),
			823 => std_logic_vector(to_unsigned(67, 8)),
			824 => std_logic_vector(to_unsigned(14, 8)),
			825 => std_logic_vector(to_unsigned(133, 8)),
			826 => std_logic_vector(to_unsigned(19, 8)),
			827 => std_logic_vector(to_unsigned(112, 8)),
			828 => std_logic_vector(to_unsigned(76, 8)),
			829 => std_logic_vector(to_unsigned(139, 8)),
			830 => std_logic_vector(to_unsigned(108, 8)),
			831 => std_logic_vector(to_unsigned(165, 8)),
			832 => std_logic_vector(to_unsigned(17, 8)),
			833 => std_logic_vector(to_unsigned(195, 8)),
			834 => std_logic_vector(to_unsigned(154, 8)),
			835 => std_logic_vector(to_unsigned(189, 8)),
			836 => std_logic_vector(to_unsigned(196, 8)),
			837 => std_logic_vector(to_unsigned(102, 8)),
			838 => std_logic_vector(to_unsigned(12, 8)),
			839 => std_logic_vector(to_unsigned(40, 8)),
			840 => std_logic_vector(to_unsigned(36, 8)),
			841 => std_logic_vector(to_unsigned(1, 8)),
			842 => std_logic_vector(to_unsigned(215, 8)),
			843 => std_logic_vector(to_unsigned(90, 8)),
			844 => std_logic_vector(to_unsigned(102, 8)),
			845 => std_logic_vector(to_unsigned(206, 8)),
			846 => std_logic_vector(to_unsigned(218, 8)),
			847 => std_logic_vector(to_unsigned(128, 8)),
			848 => std_logic_vector(to_unsigned(150, 8)),
			849 => std_logic_vector(to_unsigned(107, 8)),
			850 => std_logic_vector(to_unsigned(63, 8)),
			851 => std_logic_vector(to_unsigned(251, 8)),
			852 => std_logic_vector(to_unsigned(132, 8)),
			853 => std_logic_vector(to_unsigned(7, 8)),
			854 => std_logic_vector(to_unsigned(181, 8)),
			855 => std_logic_vector(to_unsigned(167, 8)),
			856 => std_logic_vector(to_unsigned(118, 8)),
			857 => std_logic_vector(to_unsigned(11, 8)),
			858 => std_logic_vector(to_unsigned(210, 8)),
			859 => std_logic_vector(to_unsigned(57, 8)),
			860 => std_logic_vector(to_unsigned(138, 8)),
			861 => std_logic_vector(to_unsigned(140, 8)),
			862 => std_logic_vector(to_unsigned(212, 8)),
			863 => std_logic_vector(to_unsigned(222, 8)),
			864 => std_logic_vector(to_unsigned(159, 8)),
			865 => std_logic_vector(to_unsigned(237, 8)),
			866 => std_logic_vector(to_unsigned(233, 8)),
			867 => std_logic_vector(to_unsigned(144, 8)),
			868 => std_logic_vector(to_unsigned(243, 8)),
			869 => std_logic_vector(to_unsigned(100, 8)),
			870 => std_logic_vector(to_unsigned(129, 8)),
			871 => std_logic_vector(to_unsigned(110, 8)),
			872 => std_logic_vector(to_unsigned(242, 8)),
			873 => std_logic_vector(to_unsigned(108, 8)),
			874 => std_logic_vector(to_unsigned(201, 8)),
			875 => std_logic_vector(to_unsigned(236, 8)),
			876 => std_logic_vector(to_unsigned(101, 8)),
			877 => std_logic_vector(to_unsigned(227, 8)),
			878 => std_logic_vector(to_unsigned(135, 8)),
			879 => std_logic_vector(to_unsigned(151, 8)),
			880 => std_logic_vector(to_unsigned(221, 8)),
			881 => std_logic_vector(to_unsigned(175, 8)),
			882 => std_logic_vector(to_unsigned(85, 8)),
			883 => std_logic_vector(to_unsigned(121, 8)),
			884 => std_logic_vector(to_unsigned(92, 8)),
			885 => std_logic_vector(to_unsigned(166, 8)),
			886 => std_logic_vector(to_unsigned(233, 8)),
			887 => std_logic_vector(to_unsigned(47, 8)),
			888 => std_logic_vector(to_unsigned(243, 8)),
			889 => std_logic_vector(to_unsigned(231, 8)),
			890 => std_logic_vector(to_unsigned(121, 8)),
			891 => std_logic_vector(to_unsigned(223, 8)),
			892 => std_logic_vector(to_unsigned(229, 8)),
			893 => std_logic_vector(to_unsigned(165, 8)),
			894 => std_logic_vector(to_unsigned(153, 8)),
			895 => std_logic_vector(to_unsigned(117, 8)),
			896 => std_logic_vector(to_unsigned(151, 8)),
			897 => std_logic_vector(to_unsigned(26, 8)),
			898 => std_logic_vector(to_unsigned(246, 8)),
			899 => std_logic_vector(to_unsigned(190, 8)),
			900 => std_logic_vector(to_unsigned(1, 8)),
			901 => std_logic_vector(to_unsigned(122, 8)),
			902 => std_logic_vector(to_unsigned(191, 8)),
			903 => std_logic_vector(to_unsigned(79, 8)),
			904 => std_logic_vector(to_unsigned(46, 8)),
			905 => std_logic_vector(to_unsigned(52, 8)),
			906 => std_logic_vector(to_unsigned(204, 8)),
			907 => std_logic_vector(to_unsigned(179, 8)),
			908 => std_logic_vector(to_unsigned(148, 8)),
			909 => std_logic_vector(to_unsigned(103, 8)),
			910 => std_logic_vector(to_unsigned(121, 8)),
			911 => std_logic_vector(to_unsigned(62, 8)),
			912 => std_logic_vector(to_unsigned(113, 8)),
			913 => std_logic_vector(to_unsigned(70, 8)),
			914 => std_logic_vector(to_unsigned(253, 8)),
			915 => std_logic_vector(to_unsigned(119, 8)),
			916 => std_logic_vector(to_unsigned(248, 8)),
			917 => std_logic_vector(to_unsigned(146, 8)),
			918 => std_logic_vector(to_unsigned(18, 8)),
			919 => std_logic_vector(to_unsigned(140, 8)),
			920 => std_logic_vector(to_unsigned(44, 8)),
			921 => std_logic_vector(to_unsigned(214, 8)),
			922 => std_logic_vector(to_unsigned(205, 8)),
			923 => std_logic_vector(to_unsigned(145, 8)),
			924 => std_logic_vector(to_unsigned(241, 8)),
			925 => std_logic_vector(to_unsigned(183, 8)),
			926 => std_logic_vector(to_unsigned(181, 8)),
			927 => std_logic_vector(to_unsigned(45, 8)),
			928 => std_logic_vector(to_unsigned(198, 8)),
			929 => std_logic_vector(to_unsigned(37, 8)),
			930 => std_logic_vector(to_unsigned(235, 8)),
			931 => std_logic_vector(to_unsigned(99, 8)),
			932 => std_logic_vector(to_unsigned(221, 8)),
			933 => std_logic_vector(to_unsigned(1, 8)),
			934 => std_logic_vector(to_unsigned(130, 8)),
			935 => std_logic_vector(to_unsigned(0, 8)),
			936 => std_logic_vector(to_unsigned(53, 8)),
			937 => std_logic_vector(to_unsigned(67, 8)),
			938 => std_logic_vector(to_unsigned(170, 8)),
			939 => std_logic_vector(to_unsigned(196, 8)),
			940 => std_logic_vector(to_unsigned(72, 8)),
			941 => std_logic_vector(to_unsigned(8, 8)),
			942 => std_logic_vector(to_unsigned(135, 8)),
			943 => std_logic_vector(to_unsigned(137, 8)),
			944 => std_logic_vector(to_unsigned(94, 8)),
			945 => std_logic_vector(to_unsigned(103, 8)),
			946 => std_logic_vector(to_unsigned(34, 8)),
			947 => std_logic_vector(to_unsigned(86, 8)),
			948 => std_logic_vector(to_unsigned(197, 8)),
			949 => std_logic_vector(to_unsigned(142, 8)),
			950 => std_logic_vector(to_unsigned(41, 8)),
			951 => std_logic_vector(to_unsigned(128, 8)),
			952 => std_logic_vector(to_unsigned(83, 8)),
			953 => std_logic_vector(to_unsigned(68, 8)),
			954 => std_logic_vector(to_unsigned(215, 8)),
			955 => std_logic_vector(to_unsigned(117, 8)),
			956 => std_logic_vector(to_unsigned(76, 8)),
			957 => std_logic_vector(to_unsigned(175, 8)),
			958 => std_logic_vector(to_unsigned(239, 8)),
			959 => std_logic_vector(to_unsigned(98, 8)),
			960 => std_logic_vector(to_unsigned(114, 8)),
			961 => std_logic_vector(to_unsigned(13, 8)),
			962 => std_logic_vector(to_unsigned(255, 8)),
			963 => std_logic_vector(to_unsigned(64, 8)),
			964 => std_logic_vector(to_unsigned(167, 8)),
			965 => std_logic_vector(to_unsigned(123, 8)),
			966 => std_logic_vector(to_unsigned(97, 8)),
			967 => std_logic_vector(to_unsigned(198, 8)),
			968 => std_logic_vector(to_unsigned(213, 8)),
			969 => std_logic_vector(to_unsigned(189, 8)),
			970 => std_logic_vector(to_unsigned(120, 8)),
			971 => std_logic_vector(to_unsigned(105, 8)),
			972 => std_logic_vector(to_unsigned(230, 8)),
			973 => std_logic_vector(to_unsigned(88, 8)),
			974 => std_logic_vector(to_unsigned(166, 8)),
			975 => std_logic_vector(to_unsigned(7, 8)),
			976 => std_logic_vector(to_unsigned(2, 8)),
			977 => std_logic_vector(to_unsigned(13, 8)),
			978 => std_logic_vector(to_unsigned(245, 8)),
			979 => std_logic_vector(to_unsigned(105, 8)),
			980 => std_logic_vector(to_unsigned(137, 8)),
			981 => std_logic_vector(to_unsigned(207, 8)),
			982 => std_logic_vector(to_unsigned(97, 8)),
			983 => std_logic_vector(to_unsigned(63, 8)),
			984 => std_logic_vector(to_unsigned(213, 8)),
			985 => std_logic_vector(to_unsigned(185, 8)),
			986 => std_logic_vector(to_unsigned(200, 8)),
			987 => std_logic_vector(to_unsigned(176, 8)),
			988 => std_logic_vector(to_unsigned(71, 8)),
			989 => std_logic_vector(to_unsigned(188, 8)),
			990 => std_logic_vector(to_unsigned(34, 8)),
			991 => std_logic_vector(to_unsigned(209, 8)),
			992 => std_logic_vector(to_unsigned(77, 8)),
			993 => std_logic_vector(to_unsigned(52, 8)),
			994 => std_logic_vector(to_unsigned(153, 8)),
			995 => std_logic_vector(to_unsigned(88, 8)),
			996 => std_logic_vector(to_unsigned(14, 8)),
			997 => std_logic_vector(to_unsigned(250, 8)),
			998 => std_logic_vector(to_unsigned(177, 8)),
			999 => std_logic_vector(to_unsigned(227, 8)),
			1000 => std_logic_vector(to_unsigned(204, 8)),
			1001 => std_logic_vector(to_unsigned(119, 8)),
			1002 => std_logic_vector(to_unsigned(183, 8)),
			1003 => std_logic_vector(to_unsigned(27, 8)),
			1004 => std_logic_vector(to_unsigned(219, 8)),
			1005 => std_logic_vector(to_unsigned(175, 8)),
			1006 => std_logic_vector(to_unsigned(248, 8)),
			1007 => std_logic_vector(to_unsigned(113, 8)),
			1008 => std_logic_vector(to_unsigned(50, 8)),
			1009 => std_logic_vector(to_unsigned(107, 8)),
			1010 => std_logic_vector(to_unsigned(46, 8)),
			1011 => std_logic_vector(to_unsigned(197, 8)),
			1012 => std_logic_vector(to_unsigned(16, 8)),
			1013 => std_logic_vector(to_unsigned(62, 8)),
			1014 => std_logic_vector(to_unsigned(19, 8)),
			1015 => std_logic_vector(to_unsigned(255, 8)),
			1016 => std_logic_vector(to_unsigned(177, 8)),
			1017 => std_logic_vector(to_unsigned(3, 8)),
			1018 => std_logic_vector(to_unsigned(164, 8)),
			1019 => std_logic_vector(to_unsigned(41, 8)),
			1020 => std_logic_vector(to_unsigned(167, 8)),
			1021 => std_logic_vector(to_unsigned(138, 8)),
			1022 => std_logic_vector(to_unsigned(112, 8)),
			1023 => std_logic_vector(to_unsigned(245, 8)),
			1024 => std_logic_vector(to_unsigned(16, 8)),
			1025 => std_logic_vector(to_unsigned(5, 8)),
			1026 => std_logic_vector(to_unsigned(136, 8)),
			1027 => std_logic_vector(to_unsigned(206, 8)),
			1028 => std_logic_vector(to_unsigned(82, 8)),
			1029 => std_logic_vector(to_unsigned(31, 8)),
			1030 => std_logic_vector(to_unsigned(129, 8)),
			1031 => std_logic_vector(to_unsigned(92, 8)),
			1032 => std_logic_vector(to_unsigned(155, 8)),
			1033 => std_logic_vector(to_unsigned(213, 8)),
			1034 => std_logic_vector(to_unsigned(164, 8)),
			1035 => std_logic_vector(to_unsigned(14, 8)),
			1036 => std_logic_vector(to_unsigned(233, 8)),
			1037 => std_logic_vector(to_unsigned(187, 8)),
			1038 => std_logic_vector(to_unsigned(205, 8)),
			1039 => std_logic_vector(to_unsigned(0, 8)),
			1040 => std_logic_vector(to_unsigned(192, 8)),
			1041 => std_logic_vector(to_unsigned(187, 8)),
			1042 => std_logic_vector(to_unsigned(26, 8)),
			1043 => std_logic_vector(to_unsigned(225, 8)),
			1044 => std_logic_vector(to_unsigned(4, 8)),
			1045 => std_logic_vector(to_unsigned(1, 8)),
			1046 => std_logic_vector(to_unsigned(82, 8)),
			1047 => std_logic_vector(to_unsigned(158, 8)),
			1048 => std_logic_vector(to_unsigned(248, 8)),
			1049 => std_logic_vector(to_unsigned(255, 8)),
			1050 => std_logic_vector(to_unsigned(130, 8)),
			1051 => std_logic_vector(to_unsigned(112, 8)),
			1052 => std_logic_vector(to_unsigned(176, 8)),
			1053 => std_logic_vector(to_unsigned(199, 8)),
			1054 => std_logic_vector(to_unsigned(235, 8)),
			1055 => std_logic_vector(to_unsigned(138, 8)),
			1056 => std_logic_vector(to_unsigned(28, 8)),
			1057 => std_logic_vector(to_unsigned(123, 8)),
			1058 => std_logic_vector(to_unsigned(57, 8)),
			1059 => std_logic_vector(to_unsigned(177, 8)),
			1060 => std_logic_vector(to_unsigned(233, 8)),
			1061 => std_logic_vector(to_unsigned(203, 8)),
			1062 => std_logic_vector(to_unsigned(20, 8)),
			1063 => std_logic_vector(to_unsigned(31, 8)),
			1064 => std_logic_vector(to_unsigned(112, 8)),
			1065 => std_logic_vector(to_unsigned(0, 8)),
			1066 => std_logic_vector(to_unsigned(135, 8)),
			1067 => std_logic_vector(to_unsigned(10, 8)),
			1068 => std_logic_vector(to_unsigned(202, 8)),
			1069 => std_logic_vector(to_unsigned(8, 8)),
			1070 => std_logic_vector(to_unsigned(89, 8)),
			1071 => std_logic_vector(to_unsigned(2, 8)),
			1072 => std_logic_vector(to_unsigned(40, 8)),
			1073 => std_logic_vector(to_unsigned(212, 8)),
			1074 => std_logic_vector(to_unsigned(189, 8)),
			1075 => std_logic_vector(to_unsigned(51, 8)),
			1076 => std_logic_vector(to_unsigned(39, 8)),
			1077 => std_logic_vector(to_unsigned(191, 8)),
			1078 => std_logic_vector(to_unsigned(82, 8)),
			1079 => std_logic_vector(to_unsigned(118, 8)),
			1080 => std_logic_vector(to_unsigned(237, 8)),
			1081 => std_logic_vector(to_unsigned(97, 8)),
			1082 => std_logic_vector(to_unsigned(127, 8)),
			1083 => std_logic_vector(to_unsigned(102, 8)),
			1084 => std_logic_vector(to_unsigned(71, 8)),
			1085 => std_logic_vector(to_unsigned(14, 8)),
			1086 => std_logic_vector(to_unsigned(97, 8)),
			1087 => std_logic_vector(to_unsigned(132, 8)),
			1088 => std_logic_vector(to_unsigned(17, 8)),
			1089 => std_logic_vector(to_unsigned(220, 8)),
			1090 => std_logic_vector(to_unsigned(188, 8)),
			1091 => std_logic_vector(to_unsigned(226, 8)),
			1092 => std_logic_vector(to_unsigned(3, 8)),
			1093 => std_logic_vector(to_unsigned(167, 8)),
			1094 => std_logic_vector(to_unsigned(234, 8)),
			1095 => std_logic_vector(to_unsigned(78, 8)),
			1096 => std_logic_vector(to_unsigned(2, 8)),
			1097 => std_logic_vector(to_unsigned(44, 8)),
			1098 => std_logic_vector(to_unsigned(137, 8)),
			1099 => std_logic_vector(to_unsigned(204, 8)),
			1100 => std_logic_vector(to_unsigned(211, 8)),
			1101 => std_logic_vector(to_unsigned(95, 8)),
			1102 => std_logic_vector(to_unsigned(16, 8)),
			1103 => std_logic_vector(to_unsigned(45, 8)),
			1104 => std_logic_vector(to_unsigned(218, 8)),
			1105 => std_logic_vector(to_unsigned(58, 8)),
			1106 => std_logic_vector(to_unsigned(244, 8)),
			1107 => std_logic_vector(to_unsigned(180, 8)),
			1108 => std_logic_vector(to_unsigned(110, 8)),
			1109 => std_logic_vector(to_unsigned(117, 8)),
			1110 => std_logic_vector(to_unsigned(59, 8)),
			1111 => std_logic_vector(to_unsigned(228, 8)),
			1112 => std_logic_vector(to_unsigned(32, 8)),
			1113 => std_logic_vector(to_unsigned(213, 8)),
			1114 => std_logic_vector(to_unsigned(8, 8)),
			1115 => std_logic_vector(to_unsigned(117, 8)),
			1116 => std_logic_vector(to_unsigned(181, 8)),
			1117 => std_logic_vector(to_unsigned(70, 8)),
			1118 => std_logic_vector(to_unsigned(243, 8)),
			1119 => std_logic_vector(to_unsigned(237, 8)),
			1120 => std_logic_vector(to_unsigned(68, 8)),
			1121 => std_logic_vector(to_unsigned(201, 8)),
			1122 => std_logic_vector(to_unsigned(52, 8)),
			1123 => std_logic_vector(to_unsigned(28, 8)),
			1124 => std_logic_vector(to_unsigned(243, 8)),
			1125 => std_logic_vector(to_unsigned(23, 8)),
			1126 => std_logic_vector(to_unsigned(223, 8)),
			1127 => std_logic_vector(to_unsigned(139, 8)),
			1128 => std_logic_vector(to_unsigned(250, 8)),
			1129 => std_logic_vector(to_unsigned(129, 8)),
			1130 => std_logic_vector(to_unsigned(39, 8)),
			1131 => std_logic_vector(to_unsigned(60, 8)),
			1132 => std_logic_vector(to_unsigned(13, 8)),
			1133 => std_logic_vector(to_unsigned(12, 8)),
			1134 => std_logic_vector(to_unsigned(221, 8)),
			1135 => std_logic_vector(to_unsigned(202, 8)),
			1136 => std_logic_vector(to_unsigned(241, 8)),
			1137 => std_logic_vector(to_unsigned(240, 8)),
			others => (others => '0'));
component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;
begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;
MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end process;
test : process is
begin 
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;
	assert RAM(1138) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(1138))))  severity failure;
	assert RAM(1139) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(1139))))  severity failure;
	assert RAM(1140) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(1140))))  severity failure;
	assert RAM(1141) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(1141))))  severity failure;
	assert RAM(1142) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(1142))))  severity failure;
	assert RAM(1143) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(1143))))  severity failure;
	assert RAM(1144) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(1144))))  severity failure;
	assert RAM(1145) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(1145))))  severity failure;
	assert RAM(1146) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(1146))))  severity failure;
	assert RAM(1147) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(1147))))  severity failure;
	assert RAM(1148) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(1148))))  severity failure;
	assert RAM(1149) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(1149))))  severity failure;
	assert RAM(1150) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(1150))))  severity failure;
	assert RAM(1151) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(1151))))  severity failure;
	assert RAM(1152) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(1152))))  severity failure;
	assert RAM(1153) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(1153))))  severity failure;
	assert RAM(1154) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(1154))))  severity failure;
	assert RAM(1155) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(1155))))  severity failure;
	assert RAM(1156) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(1156))))  severity failure;
	assert RAM(1157) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(1157))))  severity failure;
	assert RAM(1158) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(1158))))  severity failure;
	assert RAM(1159) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(1159))))  severity failure;
	assert RAM(1160) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(1160))))  severity failure;
	assert RAM(1161) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(1161))))  severity failure;
	assert RAM(1162) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(1162))))  severity failure;
	assert RAM(1163) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(1163))))  severity failure;
	assert RAM(1164) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(1164))))  severity failure;
	assert RAM(1165) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(1165))))  severity failure;
	assert RAM(1166) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(1166))))  severity failure;
	assert RAM(1167) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(1167))))  severity failure;
	assert RAM(1168) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(1168))))  severity failure;
	assert RAM(1169) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(1169))))  severity failure;
	assert RAM(1170) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(1170))))  severity failure;
	assert RAM(1171) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1171))))  severity failure;
	assert RAM(1172) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(1172))))  severity failure;
	assert RAM(1173) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(1173))))  severity failure;
	assert RAM(1174) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(1174))))  severity failure;
	assert RAM(1175) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(1175))))  severity failure;
	assert RAM(1176) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(1176))))  severity failure;
	assert RAM(1177) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(1177))))  severity failure;
	assert RAM(1178) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(1178))))  severity failure;
	assert RAM(1179) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(1179))))  severity failure;
	assert RAM(1180) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(1180))))  severity failure;
	assert RAM(1181) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(1181))))  severity failure;
	assert RAM(1182) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(1182))))  severity failure;
	assert RAM(1183) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(1183))))  severity failure;
	assert RAM(1184) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(1184))))  severity failure;
	assert RAM(1185) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(1185))))  severity failure;
	assert RAM(1186) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(1186))))  severity failure;
	assert RAM(1187) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1187))))  severity failure;
	assert RAM(1188) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(1188))))  severity failure;
	assert RAM(1189) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(1189))))  severity failure;
	assert RAM(1190) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(1190))))  severity failure;
	assert RAM(1191) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(1191))))  severity failure;
	assert RAM(1192) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(1192))))  severity failure;
	assert RAM(1193) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(1193))))  severity failure;
	assert RAM(1194) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(1194))))  severity failure;
	assert RAM(1195) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(1195))))  severity failure;
	assert RAM(1196) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(1196))))  severity failure;
	assert RAM(1197) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(1197))))  severity failure;
	assert RAM(1198) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(1198))))  severity failure;
	assert RAM(1199) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(1199))))  severity failure;
	assert RAM(1200) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(1200))))  severity failure;
	assert RAM(1201) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(1201))))  severity failure;
	assert RAM(1202) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(1202))))  severity failure;
	assert RAM(1203) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(1203))))  severity failure;
	assert RAM(1204) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(1204))))  severity failure;
	assert RAM(1205) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(1205))))  severity failure;
	assert RAM(1206) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(1206))))  severity failure;
	assert RAM(1207) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(1207))))  severity failure;
	assert RAM(1208) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(1208))))  severity failure;
	assert RAM(1209) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(1209))))  severity failure;
	assert RAM(1210) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(1210))))  severity failure;
	assert RAM(1211) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(1211))))  severity failure;
	assert RAM(1212) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(1212))))  severity failure;
	assert RAM(1213) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(1213))))  severity failure;
	assert RAM(1214) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(1214))))  severity failure;
	assert RAM(1215) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(1215))))  severity failure;
	assert RAM(1216) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(1216))))  severity failure;
	assert RAM(1217) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(1217))))  severity failure;
	assert RAM(1218) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1218))))  severity failure;
	assert RAM(1219) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(1219))))  severity failure;
	assert RAM(1220) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(1220))))  severity failure;
	assert RAM(1221) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(1221))))  severity failure;
	assert RAM(1222) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(1222))))  severity failure;
	assert RAM(1223) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(1223))))  severity failure;
	assert RAM(1224) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(1224))))  severity failure;
	assert RAM(1225) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(1225))))  severity failure;
	assert RAM(1226) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(1226))))  severity failure;
	assert RAM(1227) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(1227))))  severity failure;
	assert RAM(1228) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(1228))))  severity failure;
	assert RAM(1229) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(1229))))  severity failure;
	assert RAM(1230) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(1230))))  severity failure;
	assert RAM(1231) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(1231))))  severity failure;
	assert RAM(1232) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(1232))))  severity failure;
	assert RAM(1233) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(1233))))  severity failure;
	assert RAM(1234) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(1234))))  severity failure;
	assert RAM(1235) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(1235))))  severity failure;
	assert RAM(1236) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(1236))))  severity failure;
	assert RAM(1237) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(1237))))  severity failure;
	assert RAM(1238) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(1238))))  severity failure;
	assert RAM(1239) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(1239))))  severity failure;
	assert RAM(1240) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(1240))))  severity failure;
	assert RAM(1241) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(1241))))  severity failure;
	assert RAM(1242) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(1242))))  severity failure;
	assert RAM(1243) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(1243))))  severity failure;
	assert RAM(1244) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(1244))))  severity failure;
	assert RAM(1245) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(1245))))  severity failure;
	assert RAM(1246) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(1246))))  severity failure;
	assert RAM(1247) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(1247))))  severity failure;
	assert RAM(1248) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(1248))))  severity failure;
	assert RAM(1249) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(1249))))  severity failure;
	assert RAM(1250) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(1250))))  severity failure;
	assert RAM(1251) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(1251))))  severity failure;
	assert RAM(1252) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(1252))))  severity failure;
	assert RAM(1253) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(1253))))  severity failure;
	assert RAM(1254) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(1254))))  severity failure;
	assert RAM(1255) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(1255))))  severity failure;
	assert RAM(1256) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(1256))))  severity failure;
	assert RAM(1257) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(1257))))  severity failure;
	assert RAM(1258) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(1258))))  severity failure;
	assert RAM(1259) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(1259))))  severity failure;
	assert RAM(1260) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(1260))))  severity failure;
	assert RAM(1261) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(1261))))  severity failure;
	assert RAM(1262) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(1262))))  severity failure;
	assert RAM(1263) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(1263))))  severity failure;
	assert RAM(1264) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(1264))))  severity failure;
	assert RAM(1265) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(1265))))  severity failure;
	assert RAM(1266) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(1266))))  severity failure;
	assert RAM(1267) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(1267))))  severity failure;
	assert RAM(1268) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(1268))))  severity failure;
	assert RAM(1269) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(1269))))  severity failure;
	assert RAM(1270) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(1270))))  severity failure;
	assert RAM(1271) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(1271))))  severity failure;
	assert RAM(1272) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(1272))))  severity failure;
	assert RAM(1273) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(1273))))  severity failure;
	assert RAM(1274) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(1274))))  severity failure;
	assert RAM(1275) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(1275))))  severity failure;
	assert RAM(1276) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(1276))))  severity failure;
	assert RAM(1277) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(1277))))  severity failure;
	assert RAM(1278) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1278))))  severity failure;
	assert RAM(1279) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(1279))))  severity failure;
	assert RAM(1280) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(1280))))  severity failure;
	assert RAM(1281) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(1281))))  severity failure;
	assert RAM(1282) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(1282))))  severity failure;
	assert RAM(1283) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(1283))))  severity failure;
	assert RAM(1284) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(1284))))  severity failure;
	assert RAM(1285) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(1285))))  severity failure;
	assert RAM(1286) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(1286))))  severity failure;
	assert RAM(1287) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(1287))))  severity failure;
	assert RAM(1288) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(1288))))  severity failure;
	assert RAM(1289) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(1289))))  severity failure;
	assert RAM(1290) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(1290))))  severity failure;
	assert RAM(1291) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(1291))))  severity failure;
	assert RAM(1292) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(1292))))  severity failure;
	assert RAM(1293) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(1293))))  severity failure;
	assert RAM(1294) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(1294))))  severity failure;
	assert RAM(1295) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(1295))))  severity failure;
	assert RAM(1296) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(1296))))  severity failure;
	assert RAM(1297) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(1297))))  severity failure;
	assert RAM(1298) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(1298))))  severity failure;
	assert RAM(1299) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(1299))))  severity failure;
	assert RAM(1300) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1300))))  severity failure;
	assert RAM(1301) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(1301))))  severity failure;
	assert RAM(1302) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(1302))))  severity failure;
	assert RAM(1303) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(1303))))  severity failure;
	assert RAM(1304) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(1304))))  severity failure;
	assert RAM(1305) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(1305))))  severity failure;
	assert RAM(1306) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(1306))))  severity failure;
	assert RAM(1307) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(1307))))  severity failure;
	assert RAM(1308) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(1308))))  severity failure;
	assert RAM(1309) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(1309))))  severity failure;
	assert RAM(1310) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(1310))))  severity failure;
	assert RAM(1311) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(1311))))  severity failure;
	assert RAM(1312) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(1312))))  severity failure;
	assert RAM(1313) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(1313))))  severity failure;
	assert RAM(1314) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(1314))))  severity failure;
	assert RAM(1315) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(1315))))  severity failure;
	assert RAM(1316) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(1316))))  severity failure;
	assert RAM(1317) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(1317))))  severity failure;
	assert RAM(1318) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(1318))))  severity failure;
	assert RAM(1319) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(1319))))  severity failure;
	assert RAM(1320) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(1320))))  severity failure;
	assert RAM(1321) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(1321))))  severity failure;
	assert RAM(1322) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(1322))))  severity failure;
	assert RAM(1323) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(1323))))  severity failure;
	assert RAM(1324) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(1324))))  severity failure;
	assert RAM(1325) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(1325))))  severity failure;
	assert RAM(1326) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(1326))))  severity failure;
	assert RAM(1327) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(1327))))  severity failure;
	assert RAM(1328) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(1328))))  severity failure;
	assert RAM(1329) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(1329))))  severity failure;
	assert RAM(1330) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(1330))))  severity failure;
	assert RAM(1331) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(1331))))  severity failure;
	assert RAM(1332) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(1332))))  severity failure;
	assert RAM(1333) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(1333))))  severity failure;
	assert RAM(1334) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(1334))))  severity failure;
	assert RAM(1335) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(1335))))  severity failure;
	assert RAM(1336) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(1336))))  severity failure;
	assert RAM(1337) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(1337))))  severity failure;
	assert RAM(1338) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(1338))))  severity failure;
	assert RAM(1339) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(1339))))  severity failure;
	assert RAM(1340) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(1340))))  severity failure;
	assert RAM(1341) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(1341))))  severity failure;
	assert RAM(1342) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(1342))))  severity failure;
	assert RAM(1343) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(1343))))  severity failure;
	assert RAM(1344) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(1344))))  severity failure;
	assert RAM(1345) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(1345))))  severity failure;
	assert RAM(1346) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(1346))))  severity failure;
	assert RAM(1347) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(1347))))  severity failure;
	assert RAM(1348) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(1348))))  severity failure;
	assert RAM(1349) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(1349))))  severity failure;
	assert RAM(1350) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(1350))))  severity failure;
	assert RAM(1351) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(1351))))  severity failure;
	assert RAM(1352) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(1352))))  severity failure;
	assert RAM(1353) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(1353))))  severity failure;
	assert RAM(1354) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(1354))))  severity failure;
	assert RAM(1355) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(1355))))  severity failure;
	assert RAM(1356) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(1356))))  severity failure;
	assert RAM(1357) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(1357))))  severity failure;
	assert RAM(1358) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(1358))))  severity failure;
	assert RAM(1359) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(1359))))  severity failure;
	assert RAM(1360) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(1360))))  severity failure;
	assert RAM(1361) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(1361))))  severity failure;
	assert RAM(1362) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(1362))))  severity failure;
	assert RAM(1363) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(1363))))  severity failure;
	assert RAM(1364) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(1364))))  severity failure;
	assert RAM(1365) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(1365))))  severity failure;
	assert RAM(1366) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(1366))))  severity failure;
	assert RAM(1367) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(1367))))  severity failure;
	assert RAM(1368) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(1368))))  severity failure;
	assert RAM(1369) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(1369))))  severity failure;
	assert RAM(1370) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(1370))))  severity failure;
	assert RAM(1371) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(1371))))  severity failure;
	assert RAM(1372) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(1372))))  severity failure;
	assert RAM(1373) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(1373))))  severity failure;
	assert RAM(1374) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(1374))))  severity failure;
	assert RAM(1375) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(1375))))  severity failure;
	assert RAM(1376) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(1376))))  severity failure;
	assert RAM(1377) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(1377))))  severity failure;
	assert RAM(1378) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(1378))))  severity failure;
	assert RAM(1379) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(1379))))  severity failure;
	assert RAM(1380) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(1380))))  severity failure;
	assert RAM(1381) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(1381))))  severity failure;
	assert RAM(1382) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(1382))))  severity failure;
	assert RAM(1383) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(1383))))  severity failure;
	assert RAM(1384) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(1384))))  severity failure;
	assert RAM(1385) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(1385))))  severity failure;
	assert RAM(1386) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(1386))))  severity failure;
	assert RAM(1387) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(1387))))  severity failure;
	assert RAM(1388) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(1388))))  severity failure;
	assert RAM(1389) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(1389))))  severity failure;
	assert RAM(1390) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(1390))))  severity failure;
	assert RAM(1391) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(1391))))  severity failure;
	assert RAM(1392) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(1392))))  severity failure;
	assert RAM(1393) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(1393))))  severity failure;
	assert RAM(1394) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(1394))))  severity failure;
	assert RAM(1395) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(1395))))  severity failure;
	assert RAM(1396) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(1396))))  severity failure;
	assert RAM(1397) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(1397))))  severity failure;
	assert RAM(1398) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(1398))))  severity failure;
	assert RAM(1399) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(1399))))  severity failure;
	assert RAM(1400) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(1400))))  severity failure;
	assert RAM(1401) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(1401))))  severity failure;
	assert RAM(1402) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(1402))))  severity failure;
	assert RAM(1403) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(1403))))  severity failure;
	assert RAM(1404) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(1404))))  severity failure;
	assert RAM(1405) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(1405))))  severity failure;
	assert RAM(1406) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(1406))))  severity failure;
	assert RAM(1407) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(1407))))  severity failure;
	assert RAM(1408) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(1408))))  severity failure;
	assert RAM(1409) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(1409))))  severity failure;
	assert RAM(1410) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(1410))))  severity failure;
	assert RAM(1411) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(1411))))  severity failure;
	assert RAM(1412) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(1412))))  severity failure;
	assert RAM(1413) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(1413))))  severity failure;
	assert RAM(1414) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(1414))))  severity failure;
	assert RAM(1415) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(1415))))  severity failure;
	assert RAM(1416) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(1416))))  severity failure;
	assert RAM(1417) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(1417))))  severity failure;
	assert RAM(1418) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1418))))  severity failure;
	assert RAM(1419) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(1419))))  severity failure;
	assert RAM(1420) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(1420))))  severity failure;
	assert RAM(1421) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(1421))))  severity failure;
	assert RAM(1422) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(1422))))  severity failure;
	assert RAM(1423) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(1423))))  severity failure;
	assert RAM(1424) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(1424))))  severity failure;
	assert RAM(1425) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(1425))))  severity failure;
	assert RAM(1426) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(1426))))  severity failure;
	assert RAM(1427) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(1427))))  severity failure;
	assert RAM(1428) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(1428))))  severity failure;
	assert RAM(1429) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(1429))))  severity failure;
	assert RAM(1430) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(1430))))  severity failure;
	assert RAM(1431) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(1431))))  severity failure;
	assert RAM(1432) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(1432))))  severity failure;
	assert RAM(1433) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1433))))  severity failure;
	assert RAM(1434) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(1434))))  severity failure;
	assert RAM(1435) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1435))))  severity failure;
	assert RAM(1436) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(1436))))  severity failure;
	assert RAM(1437) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(1437))))  severity failure;
	assert RAM(1438) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(1438))))  severity failure;
	assert RAM(1439) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(1439))))  severity failure;
	assert RAM(1440) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(1440))))  severity failure;
	assert RAM(1441) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(1441))))  severity failure;
	assert RAM(1442) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(1442))))  severity failure;
	assert RAM(1443) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(1443))))  severity failure;
	assert RAM(1444) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(1444))))  severity failure;
	assert RAM(1445) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1445))))  severity failure;
	assert RAM(1446) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(1446))))  severity failure;
	assert RAM(1447) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(1447))))  severity failure;
	assert RAM(1448) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(1448))))  severity failure;
	assert RAM(1449) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(1449))))  severity failure;
	assert RAM(1450) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(1450))))  severity failure;
	assert RAM(1451) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(1451))))  severity failure;
	assert RAM(1452) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(1452))))  severity failure;
	assert RAM(1453) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(1453))))  severity failure;
	assert RAM(1454) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(1454))))  severity failure;
	assert RAM(1455) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(1455))))  severity failure;
	assert RAM(1456) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(1456))))  severity failure;
	assert RAM(1457) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(1457))))  severity failure;
	assert RAM(1458) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(1458))))  severity failure;
	assert RAM(1459) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(1459))))  severity failure;
	assert RAM(1460) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(1460))))  severity failure;
	assert RAM(1461) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(1461))))  severity failure;
	assert RAM(1462) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(1462))))  severity failure;
	assert RAM(1463) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(1463))))  severity failure;
	assert RAM(1464) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(1464))))  severity failure;
	assert RAM(1465) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(1465))))  severity failure;
	assert RAM(1466) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(1466))))  severity failure;
	assert RAM(1467) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(1467))))  severity failure;
	assert RAM(1468) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(1468))))  severity failure;
	assert RAM(1469) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(1469))))  severity failure;
	assert RAM(1470) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(1470))))  severity failure;
	assert RAM(1471) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(1471))))  severity failure;
	assert RAM(1472) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(1472))))  severity failure;
	assert RAM(1473) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(1473))))  severity failure;
	assert RAM(1474) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(1474))))  severity failure;
	assert RAM(1475) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(1475))))  severity failure;
	assert RAM(1476) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(1476))))  severity failure;
	assert RAM(1477) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(1477))))  severity failure;
	assert RAM(1478) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(1478))))  severity failure;
	assert RAM(1479) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(1479))))  severity failure;
	assert RAM(1480) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(1480))))  severity failure;
	assert RAM(1481) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(1481))))  severity failure;
	assert RAM(1482) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(1482))))  severity failure;
	assert RAM(1483) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(1483))))  severity failure;
	assert RAM(1484) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(1484))))  severity failure;
	assert RAM(1485) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(1485))))  severity failure;
	assert RAM(1486) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(1486))))  severity failure;
	assert RAM(1487) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(1487))))  severity failure;
	assert RAM(1488) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(1488))))  severity failure;
	assert RAM(1489) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(1489))))  severity failure;
	assert RAM(1490) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(1490))))  severity failure;
	assert RAM(1491) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(1491))))  severity failure;
	assert RAM(1492) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(1492))))  severity failure;
	assert RAM(1493) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(1493))))  severity failure;
	assert RAM(1494) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(1494))))  severity failure;
	assert RAM(1495) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(1495))))  severity failure;
	assert RAM(1496) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(1496))))  severity failure;
	assert RAM(1497) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(1497))))  severity failure;
	assert RAM(1498) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(1498))))  severity failure;
	assert RAM(1499) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(1499))))  severity failure;
	assert RAM(1500) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(1500))))  severity failure;
	assert RAM(1501) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(1501))))  severity failure;
	assert RAM(1502) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(1502))))  severity failure;
	assert RAM(1503) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(1503))))  severity failure;
	assert RAM(1504) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(1504))))  severity failure;
	assert RAM(1505) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(1505))))  severity failure;
	assert RAM(1506) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(1506))))  severity failure;
	assert RAM(1507) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(1507))))  severity failure;
	assert RAM(1508) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(1508))))  severity failure;
	assert RAM(1509) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(1509))))  severity failure;
	assert RAM(1510) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(1510))))  severity failure;
	assert RAM(1511) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(1511))))  severity failure;
	assert RAM(1512) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(1512))))  severity failure;
	assert RAM(1513) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(1513))))  severity failure;
	assert RAM(1514) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(1514))))  severity failure;
	assert RAM(1515) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(1515))))  severity failure;
	assert RAM(1516) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(1516))))  severity failure;
	assert RAM(1517) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(1517))))  severity failure;
	assert RAM(1518) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(1518))))  severity failure;
	assert RAM(1519) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(1519))))  severity failure;
	assert RAM(1520) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(1520))))  severity failure;
	assert RAM(1521) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(1521))))  severity failure;
	assert RAM(1522) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(1522))))  severity failure;
	assert RAM(1523) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(1523))))  severity failure;
	assert RAM(1524) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(1524))))  severity failure;
	assert RAM(1525) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(1525))))  severity failure;
	assert RAM(1526) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(1526))))  severity failure;
	assert RAM(1527) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(1527))))  severity failure;
	assert RAM(1528) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(1528))))  severity failure;
	assert RAM(1529) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(1529))))  severity failure;
	assert RAM(1530) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(1530))))  severity failure;
	assert RAM(1531) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(1531))))  severity failure;
	assert RAM(1532) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(1532))))  severity failure;
	assert RAM(1533) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(1533))))  severity failure;
	assert RAM(1534) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(1534))))  severity failure;
	assert RAM(1535) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(1535))))  severity failure;
	assert RAM(1536) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(1536))))  severity failure;
	assert RAM(1537) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(1537))))  severity failure;
	assert RAM(1538) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(1538))))  severity failure;
	assert RAM(1539) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(1539))))  severity failure;
	assert RAM(1540) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(1540))))  severity failure;
	assert RAM(1541) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(1541))))  severity failure;
	assert RAM(1542) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(1542))))  severity failure;
	assert RAM(1543) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(1543))))  severity failure;
	assert RAM(1544) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(1544))))  severity failure;
	assert RAM(1545) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(1545))))  severity failure;
	assert RAM(1546) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(1546))))  severity failure;
	assert RAM(1547) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(1547))))  severity failure;
	assert RAM(1548) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(1548))))  severity failure;
	assert RAM(1549) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(1549))))  severity failure;
	assert RAM(1550) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(1550))))  severity failure;
	assert RAM(1551) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(1551))))  severity failure;
	assert RAM(1552) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(1552))))  severity failure;
	assert RAM(1553) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(1553))))  severity failure;
	assert RAM(1554) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1554))))  severity failure;
	assert RAM(1555) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1555))))  severity failure;
	assert RAM(1556) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(1556))))  severity failure;
	assert RAM(1557) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(1557))))  severity failure;
	assert RAM(1558) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(1558))))  severity failure;
	assert RAM(1559) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(1559))))  severity failure;
	assert RAM(1560) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1560))))  severity failure;
	assert RAM(1561) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(1561))))  severity failure;
	assert RAM(1562) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(1562))))  severity failure;
	assert RAM(1563) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(1563))))  severity failure;
	assert RAM(1564) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(1564))))  severity failure;
	assert RAM(1565) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(1565))))  severity failure;
	assert RAM(1566) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(1566))))  severity failure;
	assert RAM(1567) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(1567))))  severity failure;
	assert RAM(1568) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(1568))))  severity failure;
	assert RAM(1569) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(1569))))  severity failure;
	assert RAM(1570) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(1570))))  severity failure;
	assert RAM(1571) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(1571))))  severity failure;
	assert RAM(1572) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(1572))))  severity failure;
	assert RAM(1573) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(1573))))  severity failure;
	assert RAM(1574) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(1574))))  severity failure;
	assert RAM(1575) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(1575))))  severity failure;
	assert RAM(1576) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(1576))))  severity failure;
	assert RAM(1577) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(1577))))  severity failure;
	assert RAM(1578) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(1578))))  severity failure;
	assert RAM(1579) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(1579))))  severity failure;
	assert RAM(1580) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(1580))))  severity failure;
	assert RAM(1581) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(1581))))  severity failure;
	assert RAM(1582) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(1582))))  severity failure;
	assert RAM(1583) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(1583))))  severity failure;
	assert RAM(1584) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(1584))))  severity failure;
	assert RAM(1585) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(1585))))  severity failure;
	assert RAM(1586) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(1586))))  severity failure;
	assert RAM(1587) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(1587))))  severity failure;
	assert RAM(1588) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(1588))))  severity failure;
	assert RAM(1589) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(1589))))  severity failure;
	assert RAM(1590) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(1590))))  severity failure;
	assert RAM(1591) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(1591))))  severity failure;
	assert RAM(1592) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(1592))))  severity failure;
	assert RAM(1593) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(1593))))  severity failure;
	assert RAM(1594) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(1594))))  severity failure;
	assert RAM(1595) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(1595))))  severity failure;
	assert RAM(1596) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(1596))))  severity failure;
	assert RAM(1597) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(1597))))  severity failure;
	assert RAM(1598) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(1598))))  severity failure;
	assert RAM(1599) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(1599))))  severity failure;
	assert RAM(1600) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(1600))))  severity failure;
	assert RAM(1601) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(1601))))  severity failure;
	assert RAM(1602) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(1602))))  severity failure;
	assert RAM(1603) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(1603))))  severity failure;
	assert RAM(1604) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(1604))))  severity failure;
	assert RAM(1605) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(1605))))  severity failure;
	assert RAM(1606) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(1606))))  severity failure;
	assert RAM(1607) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(1607))))  severity failure;
	assert RAM(1608) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(1608))))  severity failure;
	assert RAM(1609) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(1609))))  severity failure;
	assert RAM(1610) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1610))))  severity failure;
	assert RAM(1611) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(1611))))  severity failure;
	assert RAM(1612) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(1612))))  severity failure;
	assert RAM(1613) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(1613))))  severity failure;
	assert RAM(1614) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(1614))))  severity failure;
	assert RAM(1615) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(1615))))  severity failure;
	assert RAM(1616) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(1616))))  severity failure;
	assert RAM(1617) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1617))))  severity failure;
	assert RAM(1618) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(1618))))  severity failure;
	assert RAM(1619) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(1619))))  severity failure;
	assert RAM(1620) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(1620))))  severity failure;
	assert RAM(1621) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(1621))))  severity failure;
	assert RAM(1622) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(1622))))  severity failure;
	assert RAM(1623) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(1623))))  severity failure;
	assert RAM(1624) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(1624))))  severity failure;
	assert RAM(1625) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(1625))))  severity failure;
	assert RAM(1626) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(1626))))  severity failure;
	assert RAM(1627) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(1627))))  severity failure;
	assert RAM(1628) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1628))))  severity failure;
	assert RAM(1629) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(1629))))  severity failure;
	assert RAM(1630) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(1630))))  severity failure;
	assert RAM(1631) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(1631))))  severity failure;
	assert RAM(1632) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(1632))))  severity failure;
	assert RAM(1633) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(1633))))  severity failure;
	assert RAM(1634) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(1634))))  severity failure;
	assert RAM(1635) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(1635))))  severity failure;
	assert RAM(1636) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(1636))))  severity failure;
	assert RAM(1637) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(1637))))  severity failure;
	assert RAM(1638) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(1638))))  severity failure;
	assert RAM(1639) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(1639))))  severity failure;
	assert RAM(1640) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(1640))))  severity failure;
	assert RAM(1641) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(1641))))  severity failure;
	assert RAM(1642) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(1642))))  severity failure;
	assert RAM(1643) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(1643))))  severity failure;
	assert RAM(1644) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(1644))))  severity failure;
	assert RAM(1645) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(1645))))  severity failure;
	assert RAM(1646) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(1646))))  severity failure;
	assert RAM(1647) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(1647))))  severity failure;
	assert RAM(1648) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(1648))))  severity failure;
	assert RAM(1649) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(1649))))  severity failure;
	assert RAM(1650) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(1650))))  severity failure;
	assert RAM(1651) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(1651))))  severity failure;
	assert RAM(1652) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(1652))))  severity failure;
	assert RAM(1653) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(1653))))  severity failure;
	assert RAM(1654) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(1654))))  severity failure;
	assert RAM(1655) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(1655))))  severity failure;
	assert RAM(1656) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(1656))))  severity failure;
	assert RAM(1657) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(1657))))  severity failure;
	assert RAM(1658) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(1658))))  severity failure;
	assert RAM(1659) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(1659))))  severity failure;
	assert RAM(1660) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(1660))))  severity failure;
	assert RAM(1661) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(1661))))  severity failure;
	assert RAM(1662) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(1662))))  severity failure;
	assert RAM(1663) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(1663))))  severity failure;
	assert RAM(1664) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(1664))))  severity failure;
	assert RAM(1665) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(1665))))  severity failure;
	assert RAM(1666) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(1666))))  severity failure;
	assert RAM(1667) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(1667))))  severity failure;
	assert RAM(1668) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(1668))))  severity failure;
	assert RAM(1669) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(1669))))  severity failure;
	assert RAM(1670) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(1670))))  severity failure;
	assert RAM(1671) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(1671))))  severity failure;
	assert RAM(1672) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(1672))))  severity failure;
	assert RAM(1673) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(1673))))  severity failure;
	assert RAM(1674) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(1674))))  severity failure;
	assert RAM(1675) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(1675))))  severity failure;
	assert RAM(1676) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(1676))))  severity failure;
	assert RAM(1677) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(1677))))  severity failure;
	assert RAM(1678) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(1678))))  severity failure;
	assert RAM(1679) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(1679))))  severity failure;
	assert RAM(1680) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(1680))))  severity failure;
	assert RAM(1681) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(1681))))  severity failure;
	assert RAM(1682) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(1682))))  severity failure;
	assert RAM(1683) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(1683))))  severity failure;
	assert RAM(1684) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(1684))))  severity failure;
	assert RAM(1685) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(1685))))  severity failure;
	assert RAM(1686) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(1686))))  severity failure;
	assert RAM(1687) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(1687))))  severity failure;
	assert RAM(1688) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(1688))))  severity failure;
	assert RAM(1689) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(1689))))  severity failure;
	assert RAM(1690) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(1690))))  severity failure;
	assert RAM(1691) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(1691))))  severity failure;
	assert RAM(1692) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(1692))))  severity failure;
	assert RAM(1693) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(1693))))  severity failure;
	assert RAM(1694) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(1694))))  severity failure;
	assert RAM(1695) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(1695))))  severity failure;
	assert RAM(1696) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(1696))))  severity failure;
	assert RAM(1697) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(1697))))  severity failure;
	assert RAM(1698) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(1698))))  severity failure;
	assert RAM(1699) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(1699))))  severity failure;
	assert RAM(1700) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(1700))))  severity failure;
	assert RAM(1701) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(1701))))  severity failure;
	assert RAM(1702) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(1702))))  severity failure;
	assert RAM(1703) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(1703))))  severity failure;
	assert RAM(1704) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(1704))))  severity failure;
	assert RAM(1705) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(1705))))  severity failure;
	assert RAM(1706) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(1706))))  severity failure;
	assert RAM(1707) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(1707))))  severity failure;
	assert RAM(1708) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(1708))))  severity failure;
	assert RAM(1709) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(1709))))  severity failure;
	assert RAM(1710) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(1710))))  severity failure;
	assert RAM(1711) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(1711))))  severity failure;
	assert RAM(1712) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(1712))))  severity failure;
	assert RAM(1713) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(1713))))  severity failure;
	assert RAM(1714) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(1714))))  severity failure;
	assert RAM(1715) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(1715))))  severity failure;
	assert RAM(1716) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(1716))))  severity failure;
	assert RAM(1717) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(1717))))  severity failure;
	assert RAM(1718) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(1718))))  severity failure;
	assert RAM(1719) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(1719))))  severity failure;
	assert RAM(1720) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(1720))))  severity failure;
	assert RAM(1721) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(1721))))  severity failure;
	assert RAM(1722) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(1722))))  severity failure;
	assert RAM(1723) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(1723))))  severity failure;
	assert RAM(1724) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(1724))))  severity failure;
	assert RAM(1725) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(1725))))  severity failure;
	assert RAM(1726) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(1726))))  severity failure;
	assert RAM(1727) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(1727))))  severity failure;
	assert RAM(1728) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(1728))))  severity failure;
	assert RAM(1729) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(1729))))  severity failure;
	assert RAM(1730) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(1730))))  severity failure;
	assert RAM(1731) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(1731))))  severity failure;
	assert RAM(1732) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(1732))))  severity failure;
	assert RAM(1733) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(1733))))  severity failure;
	assert RAM(1734) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(1734))))  severity failure;
	assert RAM(1735) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(1735))))  severity failure;
	assert RAM(1736) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(1736))))  severity failure;
	assert RAM(1737) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(1737))))  severity failure;
	assert RAM(1738) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(1738))))  severity failure;
	assert RAM(1739) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(1739))))  severity failure;
	assert RAM(1740) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(1740))))  severity failure;
	assert RAM(1741) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(1741))))  severity failure;
	assert RAM(1742) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(1742))))  severity failure;
	assert RAM(1743) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(1743))))  severity failure;
	assert RAM(1744) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(1744))))  severity failure;
	assert RAM(1745) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(1745))))  severity failure;
	assert RAM(1746) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(1746))))  severity failure;
	assert RAM(1747) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(1747))))  severity failure;
	assert RAM(1748) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1748))))  severity failure;
	assert RAM(1749) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(1749))))  severity failure;
	assert RAM(1750) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(1750))))  severity failure;
	assert RAM(1751) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(1751))))  severity failure;
	assert RAM(1752) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(1752))))  severity failure;
	assert RAM(1753) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(1753))))  severity failure;
	assert RAM(1754) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(1754))))  severity failure;
	assert RAM(1755) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(1755))))  severity failure;
	assert RAM(1756) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(1756))))  severity failure;
	assert RAM(1757) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(1757))))  severity failure;
	assert RAM(1758) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(1758))))  severity failure;
	assert RAM(1759) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(1759))))  severity failure;
	assert RAM(1760) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(1760))))  severity failure;
	assert RAM(1761) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(1761))))  severity failure;
	assert RAM(1762) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(1762))))  severity failure;
	assert RAM(1763) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(1763))))  severity failure;
	assert RAM(1764) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(1764))))  severity failure;
	assert RAM(1765) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(1765))))  severity failure;
	assert RAM(1766) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(1766))))  severity failure;
	assert RAM(1767) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(1767))))  severity failure;
	assert RAM(1768) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(1768))))  severity failure;
	assert RAM(1769) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(1769))))  severity failure;
	assert RAM(1770) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(1770))))  severity failure;
	assert RAM(1771) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(1771))))  severity failure;
	assert RAM(1772) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(1772))))  severity failure;
	assert RAM(1773) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(1773))))  severity failure;
	assert RAM(1774) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(1774))))  severity failure;
	assert RAM(1775) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(1775))))  severity failure;
	assert RAM(1776) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(1776))))  severity failure;
	assert RAM(1777) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(1777))))  severity failure;
	assert RAM(1778) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(1778))))  severity failure;
	assert RAM(1779) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(1779))))  severity failure;
	assert RAM(1780) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(1780))))  severity failure;
	assert RAM(1781) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(1781))))  severity failure;
	assert RAM(1782) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(1782))))  severity failure;
	assert RAM(1783) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(1783))))  severity failure;
	assert RAM(1784) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(1784))))  severity failure;
	assert RAM(1785) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(1785))))  severity failure;
	assert RAM(1786) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(1786))))  severity failure;
	assert RAM(1787) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(1787))))  severity failure;
	assert RAM(1788) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(1788))))  severity failure;
	assert RAM(1789) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(1789))))  severity failure;
	assert RAM(1790) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(1790))))  severity failure;
	assert RAM(1791) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(1791))))  severity failure;
	assert RAM(1792) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(1792))))  severity failure;
	assert RAM(1793) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(1793))))  severity failure;
	assert RAM(1794) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1794))))  severity failure;
	assert RAM(1795) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(1795))))  severity failure;
	assert RAM(1796) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(1796))))  severity failure;
	assert RAM(1797) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(1797))))  severity failure;
	assert RAM(1798) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(1798))))  severity failure;
	assert RAM(1799) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(1799))))  severity failure;
	assert RAM(1800) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(1800))))  severity failure;
	assert RAM(1801) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(1801))))  severity failure;
	assert RAM(1802) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(1802))))  severity failure;
	assert RAM(1803) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(1803))))  severity failure;
	assert RAM(1804) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(1804))))  severity failure;
	assert RAM(1805) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(1805))))  severity failure;
	assert RAM(1806) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(1806))))  severity failure;
	assert RAM(1807) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(1807))))  severity failure;
	assert RAM(1808) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(1808))))  severity failure;
	assert RAM(1809) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(1809))))  severity failure;
	assert RAM(1810) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1810))))  severity failure;
	assert RAM(1811) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(1811))))  severity failure;
	assert RAM(1812) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(1812))))  severity failure;
	assert RAM(1813) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(1813))))  severity failure;
	assert RAM(1814) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(1814))))  severity failure;
	assert RAM(1815) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(1815))))  severity failure;
	assert RAM(1816) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(1816))))  severity failure;
	assert RAM(1817) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(1817))))  severity failure;
	assert RAM(1818) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(1818))))  severity failure;
	assert RAM(1819) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(1819))))  severity failure;
	assert RAM(1820) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(1820))))  severity failure;
	assert RAM(1821) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(1821))))  severity failure;
	assert RAM(1822) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(1822))))  severity failure;
	assert RAM(1823) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(1823))))  severity failure;
	assert RAM(1824) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(1824))))  severity failure;
	assert RAM(1825) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(1825))))  severity failure;
	assert RAM(1826) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(1826))))  severity failure;
	assert RAM(1827) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(1827))))  severity failure;
	assert RAM(1828) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(1828))))  severity failure;
	assert RAM(1829) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(1829))))  severity failure;
	assert RAM(1830) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(1830))))  severity failure;
	assert RAM(1831) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(1831))))  severity failure;
	assert RAM(1832) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(1832))))  severity failure;
	assert RAM(1833) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(1833))))  severity failure;
	assert RAM(1834) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(1834))))  severity failure;
	assert RAM(1835) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(1835))))  severity failure;
	assert RAM(1836) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(1836))))  severity failure;
	assert RAM(1837) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(1837))))  severity failure;
	assert RAM(1838) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(1838))))  severity failure;
	assert RAM(1839) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(1839))))  severity failure;
	assert RAM(1840) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(1840))))  severity failure;
	assert RAM(1841) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(1841))))  severity failure;
	assert RAM(1842) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(1842))))  severity failure;
	assert RAM(1843) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(1843))))  severity failure;
	assert RAM(1844) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(1844))))  severity failure;
	assert RAM(1845) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(1845))))  severity failure;
	assert RAM(1846) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(1846))))  severity failure;
	assert RAM(1847) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(1847))))  severity failure;
	assert RAM(1848) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(1848))))  severity failure;
	assert RAM(1849) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(1849))))  severity failure;
	assert RAM(1850) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(1850))))  severity failure;
	assert RAM(1851) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(1851))))  severity failure;
	assert RAM(1852) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(1852))))  severity failure;
	assert RAM(1853) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(1853))))  severity failure;
	assert RAM(1854) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(1854))))  severity failure;
	assert RAM(1855) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(1855))))  severity failure;
	assert RAM(1856) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(1856))))  severity failure;
	assert RAM(1857) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(1857))))  severity failure;
	assert RAM(1858) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(1858))))  severity failure;
	assert RAM(1859) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(1859))))  severity failure;
	assert RAM(1860) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(1860))))  severity failure;
	assert RAM(1861) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(1861))))  severity failure;
	assert RAM(1862) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(1862))))  severity failure;
	assert RAM(1863) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(1863))))  severity failure;
	assert RAM(1864) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(1864))))  severity failure;
	assert RAM(1865) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(1865))))  severity failure;
	assert RAM(1866) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(1866))))  severity failure;
	assert RAM(1867) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(1867))))  severity failure;
	assert RAM(1868) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(1868))))  severity failure;
	assert RAM(1869) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(1869))))  severity failure;
	assert RAM(1870) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(1870))))  severity failure;
	assert RAM(1871) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(1871))))  severity failure;
	assert RAM(1872) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(1872))))  severity failure;
	assert RAM(1873) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(1873))))  severity failure;
	assert RAM(1874) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(1874))))  severity failure;
	assert RAM(1875) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(1875))))  severity failure;
	assert RAM(1876) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(1876))))  severity failure;
	assert RAM(1877) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(1877))))  severity failure;
	assert RAM(1878) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(1878))))  severity failure;
	assert RAM(1879) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(1879))))  severity failure;
	assert RAM(1880) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(1880))))  severity failure;
	assert RAM(1881) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(1881))))  severity failure;
	assert RAM(1882) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(1882))))  severity failure;
	assert RAM(1883) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(1883))))  severity failure;
	assert RAM(1884) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(1884))))  severity failure;
	assert RAM(1885) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(1885))))  severity failure;
	assert RAM(1886) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(1886))))  severity failure;
	assert RAM(1887) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(1887))))  severity failure;
	assert RAM(1888) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(1888))))  severity failure;
	assert RAM(1889) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(1889))))  severity failure;
	assert RAM(1890) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(1890))))  severity failure;
	assert RAM(1891) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(1891))))  severity failure;
	assert RAM(1892) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(1892))))  severity failure;
	assert RAM(1893) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(1893))))  severity failure;
	assert RAM(1894) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(1894))))  severity failure;
	assert RAM(1895) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(1895))))  severity failure;
	assert RAM(1896) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(1896))))  severity failure;
	assert RAM(1897) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(1897))))  severity failure;
	assert RAM(1898) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(1898))))  severity failure;
	assert RAM(1899) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(1899))))  severity failure;
	assert RAM(1900) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(1900))))  severity failure;
	assert RAM(1901) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(1901))))  severity failure;
	assert RAM(1902) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(1902))))  severity failure;
	assert RAM(1903) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(1903))))  severity failure;
	assert RAM(1904) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(1904))))  severity failure;
	assert RAM(1905) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(1905))))  severity failure;
	assert RAM(1906) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(1906))))  severity failure;
	assert RAM(1907) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(1907))))  severity failure;
	assert RAM(1908) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(1908))))  severity failure;
	assert RAM(1909) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(1909))))  severity failure;
	assert RAM(1910) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(1910))))  severity failure;
	assert RAM(1911) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(1911))))  severity failure;
	assert RAM(1912) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(1912))))  severity failure;
	assert RAM(1913) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(1913))))  severity failure;
	assert RAM(1914) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(1914))))  severity failure;
	assert RAM(1915) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(1915))))  severity failure;
	assert RAM(1916) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(1916))))  severity failure;
	assert RAM(1917) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(1917))))  severity failure;
	assert RAM(1918) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(1918))))  severity failure;
	assert RAM(1919) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(1919))))  severity failure;
	assert RAM(1920) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(1920))))  severity failure;
	assert RAM(1921) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(1921))))  severity failure;
	assert RAM(1922) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(1922))))  severity failure;
	assert RAM(1923) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(1923))))  severity failure;
	assert RAM(1924) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(1924))))  severity failure;
	assert RAM(1925) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(1925))))  severity failure;
	assert RAM(1926) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(1926))))  severity failure;
	assert RAM(1927) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(1927))))  severity failure;
	assert RAM(1928) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(1928))))  severity failure;
	assert RAM(1929) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(1929))))  severity failure;
	assert RAM(1930) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(1930))))  severity failure;
	assert RAM(1931) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(1931))))  severity failure;
	assert RAM(1932) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(1932))))  severity failure;
	assert RAM(1933) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(1933))))  severity failure;
	assert RAM(1934) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(1934))))  severity failure;
	assert RAM(1935) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(1935))))  severity failure;
	assert RAM(1936) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(1936))))  severity failure;
	assert RAM(1937) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(1937))))  severity failure;
	assert RAM(1938) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(1938))))  severity failure;
	assert RAM(1939) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(1939))))  severity failure;
	assert RAM(1940) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(1940))))  severity failure;
	assert RAM(1941) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(1941))))  severity failure;
	assert RAM(1942) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(1942))))  severity failure;
	assert RAM(1943) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(1943))))  severity failure;
	assert RAM(1944) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(1944))))  severity failure;
	assert RAM(1945) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(1945))))  severity failure;
	assert RAM(1946) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(1946))))  severity failure;
	assert RAM(1947) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(1947))))  severity failure;
	assert RAM(1948) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(1948))))  severity failure;
	assert RAM(1949) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(1949))))  severity failure;
	assert RAM(1950) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(1950))))  severity failure;
	assert RAM(1951) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(1951))))  severity failure;
	assert RAM(1952) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(1952))))  severity failure;
	assert RAM(1953) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(1953))))  severity failure;
	assert RAM(1954) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(1954))))  severity failure;
	assert RAM(1955) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(1955))))  severity failure;
	assert RAM(1956) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(1956))))  severity failure;
	assert RAM(1957) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(1957))))  severity failure;
	assert RAM(1958) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(1958))))  severity failure;
	assert RAM(1959) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(1959))))  severity failure;
	assert RAM(1960) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(1960))))  severity failure;
	assert RAM(1961) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(1961))))  severity failure;
	assert RAM(1962) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(1962))))  severity failure;
	assert RAM(1963) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(1963))))  severity failure;
	assert RAM(1964) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(1964))))  severity failure;
	assert RAM(1965) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(1965))))  severity failure;
	assert RAM(1966) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(1966))))  severity failure;
	assert RAM(1967) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(1967))))  severity failure;
	assert RAM(1968) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(1968))))  severity failure;
	assert RAM(1969) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(1969))))  severity failure;
	assert RAM(1970) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(1970))))  severity failure;
	assert RAM(1971) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(1971))))  severity failure;
	assert RAM(1972) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(1972))))  severity failure;
	assert RAM(1973) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(1973))))  severity failure;
	assert RAM(1974) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(1974))))  severity failure;
	assert RAM(1975) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(1975))))  severity failure;
	assert RAM(1976) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(1976))))  severity failure;
	assert RAM(1977) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(1977))))  severity failure;
	assert RAM(1978) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(1978))))  severity failure;
	assert RAM(1979) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(1979))))  severity failure;
	assert RAM(1980) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(1980))))  severity failure;
	assert RAM(1981) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(1981))))  severity failure;
	assert RAM(1982) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(1982))))  severity failure;
	assert RAM(1983) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(1983))))  severity failure;
	assert RAM(1984) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(1984))))  severity failure;
	assert RAM(1985) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(1985))))  severity failure;
	assert RAM(1986) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(1986))))  severity failure;
	assert RAM(1987) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(1987))))  severity failure;
	assert RAM(1988) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(1988))))  severity failure;
	assert RAM(1989) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(1989))))  severity failure;
	assert RAM(1990) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(1990))))  severity failure;
	assert RAM(1991) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(1991))))  severity failure;
	assert RAM(1992) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(1992))))  severity failure;
	assert RAM(1993) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(1993))))  severity failure;
	assert RAM(1994) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(1994))))  severity failure;
	assert RAM(1995) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(1995))))  severity failure;
	assert RAM(1996) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(1996))))  severity failure;
	assert RAM(1997) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(1997))))  severity failure;
	assert RAM(1998) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(1998))))  severity failure;
	assert RAM(1999) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(1999))))  severity failure;
	assert RAM(2000) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(2000))))  severity failure;
	assert RAM(2001) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(2001))))  severity failure;
	assert RAM(2002) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2002))))  severity failure;
	assert RAM(2003) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(2003))))  severity failure;
	assert RAM(2004) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(2004))))  severity failure;
	assert RAM(2005) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(2005))))  severity failure;
	assert RAM(2006) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2006))))  severity failure;
	assert RAM(2007) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(2007))))  severity failure;
	assert RAM(2008) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(2008))))  severity failure;
	assert RAM(2009) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(2009))))  severity failure;
	assert RAM(2010) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(2010))))  severity failure;
	assert RAM(2011) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(2011))))  severity failure;
	assert RAM(2012) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(2012))))  severity failure;
	assert RAM(2013) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(2013))))  severity failure;
	assert RAM(2014) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(2014))))  severity failure;
	assert RAM(2015) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2015))))  severity failure;
	assert RAM(2016) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(2016))))  severity failure;
	assert RAM(2017) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(2017))))  severity failure;
	assert RAM(2018) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(2018))))  severity failure;
	assert RAM(2019) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2019))))  severity failure;
	assert RAM(2020) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(2020))))  severity failure;
	assert RAM(2021) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(2021))))  severity failure;
	assert RAM(2022) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2022))))  severity failure;
	assert RAM(2023) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(2023))))  severity failure;
	assert RAM(2024) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(2024))))  severity failure;
	assert RAM(2025) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(2025))))  severity failure;
	assert RAM(2026) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2026))))  severity failure;
	assert RAM(2027) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2027))))  severity failure;
	assert RAM(2028) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2028))))  severity failure;
	assert RAM(2029) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(2029))))  severity failure;
	assert RAM(2030) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(2030))))  severity failure;
	assert RAM(2031) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(2031))))  severity failure;
	assert RAM(2032) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2032))))  severity failure;
	assert RAM(2033) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2033))))  severity failure;
	assert RAM(2034) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(2034))))  severity failure;
	assert RAM(2035) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(2035))))  severity failure;
	assert RAM(2036) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(2036))))  severity failure;
	assert RAM(2037) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(2037))))  severity failure;
	assert RAM(2038) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(2038))))  severity failure;
	assert RAM(2039) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(2039))))  severity failure;
	assert RAM(2040) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(2040))))  severity failure;
	assert RAM(2041) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(2041))))  severity failure;
	assert RAM(2042) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(2042))))  severity failure;
	assert RAM(2043) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(2043))))  severity failure;
	assert RAM(2044) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(2044))))  severity failure;
	assert RAM(2045) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(2045))))  severity failure;
	assert RAM(2046) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2046))))  severity failure;
	assert RAM(2047) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(2047))))  severity failure;
	assert RAM(2048) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(2048))))  severity failure;
	assert RAM(2049) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(2049))))  severity failure;
	assert RAM(2050) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(2050))))  severity failure;
	assert RAM(2051) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(2051))))  severity failure;
	assert RAM(2052) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2052))))  severity failure;
	assert RAM(2053) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2053))))  severity failure;
	assert RAM(2054) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(2054))))  severity failure;
	assert RAM(2055) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(2055))))  severity failure;
	assert RAM(2056) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(2056))))  severity failure;
	assert RAM(2057) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(2057))))  severity failure;
	assert RAM(2058) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2058))))  severity failure;
	assert RAM(2059) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2059))))  severity failure;
	assert RAM(2060) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(2060))))  severity failure;
	assert RAM(2061) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2061))))  severity failure;
	assert RAM(2062) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(2062))))  severity failure;
	assert RAM(2063) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(2063))))  severity failure;
	assert RAM(2064) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(2064))))  severity failure;
	assert RAM(2065) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(2065))))  severity failure;
	assert RAM(2066) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(2066))))  severity failure;
	assert RAM(2067) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(2067))))  severity failure;
	assert RAM(2068) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(2068))))  severity failure;
	assert RAM(2069) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(2069))))  severity failure;
	assert RAM(2070) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(2070))))  severity failure;
	assert RAM(2071) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(2071))))  severity failure;
	assert RAM(2072) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(2072))))  severity failure;
	assert RAM(2073) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(2073))))  severity failure;
	assert RAM(2074) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(2074))))  severity failure;
	assert RAM(2075) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(2075))))  severity failure;
	assert RAM(2076) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(2076))))  severity failure;
	assert RAM(2077) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2077))))  severity failure;
	assert RAM(2078) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(2078))))  severity failure;
	assert RAM(2079) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(2079))))  severity failure;
	assert RAM(2080) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(2080))))  severity failure;
	assert RAM(2081) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(2081))))  severity failure;
	assert RAM(2082) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(2082))))  severity failure;
	assert RAM(2083) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(2083))))  severity failure;
	assert RAM(2084) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(2084))))  severity failure;
	assert RAM(2085) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(2085))))  severity failure;
	assert RAM(2086) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(2086))))  severity failure;
	assert RAM(2087) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(2087))))  severity failure;
	assert RAM(2088) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(2088))))  severity failure;
	assert RAM(2089) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(2089))))  severity failure;
	assert RAM(2090) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(2090))))  severity failure;
	assert RAM(2091) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(2091))))  severity failure;
	assert RAM(2092) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(2092))))  severity failure;
	assert RAM(2093) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(2093))))  severity failure;
	assert RAM(2094) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(2094))))  severity failure;
	assert RAM(2095) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2095))))  severity failure;
	assert RAM(2096) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(2096))))  severity failure;
	assert RAM(2097) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(2097))))  severity failure;
	assert RAM(2098) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2098))))  severity failure;
	assert RAM(2099) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(2099))))  severity failure;
	assert RAM(2100) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(2100))))  severity failure;
	assert RAM(2101) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2101))))  severity failure;
	assert RAM(2102) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(2102))))  severity failure;
	assert RAM(2103) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(2103))))  severity failure;
	assert RAM(2104) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(2104))))  severity failure;
	assert RAM(2105) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(2105))))  severity failure;
	assert RAM(2106) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(2106))))  severity failure;
	assert RAM(2107) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(2107))))  severity failure;
	assert RAM(2108) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(2108))))  severity failure;
	assert RAM(2109) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(2109))))  severity failure;
	assert RAM(2110) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(2110))))  severity failure;
	assert RAM(2111) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(2111))))  severity failure;
	assert RAM(2112) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(2112))))  severity failure;
	assert RAM(2113) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(2113))))  severity failure;
	assert RAM(2114) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2114))))  severity failure;
	assert RAM(2115) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(2115))))  severity failure;
	assert RAM(2116) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(2116))))  severity failure;
	assert RAM(2117) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(2117))))  severity failure;
	assert RAM(2118) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(2118))))  severity failure;
	assert RAM(2119) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(2119))))  severity failure;
	assert RAM(2120) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(2120))))  severity failure;
	assert RAM(2121) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(2121))))  severity failure;
	assert RAM(2122) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2122))))  severity failure;
	assert RAM(2123) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(2123))))  severity failure;
	assert RAM(2124) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(2124))))  severity failure;
	assert RAM(2125) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(2125))))  severity failure;
	assert RAM(2126) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(2126))))  severity failure;
	assert RAM(2127) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2127))))  severity failure;
	assert RAM(2128) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(2128))))  severity failure;
	assert RAM(2129) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(2129))))  severity failure;
	assert RAM(2130) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(2130))))  severity failure;
	assert RAM(2131) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(2131))))  severity failure;
	assert RAM(2132) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2132))))  severity failure;
	assert RAM(2133) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(2133))))  severity failure;
	assert RAM(2134) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(2134))))  severity failure;
	assert RAM(2135) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(2135))))  severity failure;
	assert RAM(2136) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(2136))))  severity failure;
	assert RAM(2137) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(2137))))  severity failure;
	assert RAM(2138) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2138))))  severity failure;
	assert RAM(2139) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2139))))  severity failure;
	assert RAM(2140) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(2140))))  severity failure;
	assert RAM(2141) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(2141))))  severity failure;
	assert RAM(2142) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2142))))  severity failure;
	assert RAM(2143) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(2143))))  severity failure;
	assert RAM(2144) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(2144))))  severity failure;
	assert RAM(2145) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(2145))))  severity failure;
	assert RAM(2146) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(2146))))  severity failure;
	assert RAM(2147) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(2147))))  severity failure;
	assert RAM(2148) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(2148))))  severity failure;
	assert RAM(2149) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(2149))))  severity failure;
	assert RAM(2150) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(2150))))  severity failure;
	assert RAM(2151) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2151))))  severity failure;
	assert RAM(2152) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(2152))))  severity failure;
	assert RAM(2153) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(2153))))  severity failure;
	assert RAM(2154) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(2154))))  severity failure;
	assert RAM(2155) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(2155))))  severity failure;
	assert RAM(2156) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(2156))))  severity failure;
	assert RAM(2157) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(2157))))  severity failure;
	assert RAM(2158) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2158))))  severity failure;
	assert RAM(2159) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2159))))  severity failure;
	assert RAM(2160) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(2160))))  severity failure;
	assert RAM(2161) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(2161))))  severity failure;
	assert RAM(2162) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(2162))))  severity failure;
	assert RAM(2163) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(2163))))  severity failure;
	assert RAM(2164) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(2164))))  severity failure;
	assert RAM(2165) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(2165))))  severity failure;
	assert RAM(2166) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2166))))  severity failure;
	assert RAM(2167) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(2167))))  severity failure;
	assert RAM(2168) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(2168))))  severity failure;
	assert RAM(2169) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(2169))))  severity failure;
	assert RAM(2170) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(2170))))  severity failure;
	assert RAM(2171) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2171))))  severity failure;
	assert RAM(2172) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2172))))  severity failure;
	assert RAM(2173) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(2173))))  severity failure;
	assert RAM(2174) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2174))))  severity failure;
	assert RAM(2175) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(2175))))  severity failure;
	assert RAM(2176) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(2176))))  severity failure;
	assert RAM(2177) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(2177))))  severity failure;
	assert RAM(2178) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2178))))  severity failure;
	assert RAM(2179) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(2179))))  severity failure;
	assert RAM(2180) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(2180))))  severity failure;
	assert RAM(2181) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(2181))))  severity failure;
	assert RAM(2182) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(2182))))  severity failure;
	assert RAM(2183) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(2183))))  severity failure;
	assert RAM(2184) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2184))))  severity failure;
	assert RAM(2185) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2185))))  severity failure;
	assert RAM(2186) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(2186))))  severity failure;
	assert RAM(2187) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2187))))  severity failure;
	assert RAM(2188) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(2188))))  severity failure;
	assert RAM(2189) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(2189))))  severity failure;
	assert RAM(2190) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(2190))))  severity failure;
	assert RAM(2191) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(2191))))  severity failure;
	assert RAM(2192) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(2192))))  severity failure;
	assert RAM(2193) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2193))))  severity failure;
	assert RAM(2194) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(2194))))  severity failure;
	assert RAM(2195) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(2195))))  severity failure;
	assert RAM(2196) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2196))))  severity failure;
	assert RAM(2197) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(2197))))  severity failure;
	assert RAM(2198) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(2198))))  severity failure;
	assert RAM(2199) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(2199))))  severity failure;
	assert RAM(2200) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2200))))  severity failure;
	assert RAM(2201) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(2201))))  severity failure;
	assert RAM(2202) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(2202))))  severity failure;
	assert RAM(2203) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(2203))))  severity failure;
	assert RAM(2204) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2204))))  severity failure;
	assert RAM(2205) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2205))))  severity failure;
	assert RAM(2206) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(2206))))  severity failure;
	assert RAM(2207) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(2207))))  severity failure;
	assert RAM(2208) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(2208))))  severity failure;
	assert RAM(2209) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(2209))))  severity failure;
	assert RAM(2210) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(2210))))  severity failure;
	assert RAM(2211) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(2211))))  severity failure;
	assert RAM(2212) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(2212))))  severity failure;
	assert RAM(2213) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(2213))))  severity failure;
	assert RAM(2214) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(2214))))  severity failure;
	assert RAM(2215) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(2215))))  severity failure;
	assert RAM(2216) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(2216))))  severity failure;
	assert RAM(2217) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(2217))))  severity failure;
	assert RAM(2218) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(2218))))  severity failure;
	assert RAM(2219) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2219))))  severity failure;
	assert RAM(2220) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(2220))))  severity failure;
	assert RAM(2221) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2221))))  severity failure;
	assert RAM(2222) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(2222))))  severity failure;
	assert RAM(2223) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(2223))))  severity failure;
	assert RAM(2224) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(2224))))  severity failure;
	assert RAM(2225) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(2225))))  severity failure;
	assert RAM(2226) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(2226))))  severity failure;
	assert RAM(2227) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(2227))))  severity failure;
	assert RAM(2228) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(2228))))  severity failure;
	assert RAM(2229) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(2229))))  severity failure;
	assert RAM(2230) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(2230))))  severity failure;
	assert RAM(2231) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(2231))))  severity failure;
	assert RAM(2232) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(2232))))  severity failure;
	assert RAM(2233) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(2233))))  severity failure;
	assert RAM(2234) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(2234))))  severity failure;
	assert RAM(2235) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(2235))))  severity failure;
	assert RAM(2236) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(2236))))  severity failure;
	assert RAM(2237) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(2237))))  severity failure;
	assert RAM(2238) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(2238))))  severity failure;
	assert RAM(2239) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(2239))))  severity failure;
	assert RAM(2240) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(2240))))  severity failure;
	assert RAM(2241) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(2241))))  severity failure;
	assert RAM(2242) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(2242))))  severity failure;
	assert RAM(2243) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(2243))))  severity failure;
	assert RAM(2244) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(2244))))  severity failure;
	assert RAM(2245) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(2245))))  severity failure;
	assert RAM(2246) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(2246))))  severity failure;
	assert RAM(2247) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(2247))))  severity failure;
	assert RAM(2248) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(2248))))  severity failure;
	assert RAM(2249) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(2249))))  severity failure;
	assert RAM(2250) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2250))))  severity failure;
	assert RAM(2251) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(2251))))  severity failure;
	assert RAM(2252) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(2252))))  severity failure;
	assert RAM(2253) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(2253))))  severity failure;
	assert RAM(2254) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(2254))))  severity failure;
	assert RAM(2255) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(2255))))  severity failure;
	assert RAM(2256) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(2256))))  severity failure;
	assert RAM(2257) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(2257))))  severity failure;
	assert RAM(2258) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(2258))))  severity failure;
	assert RAM(2259) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(2259))))  severity failure;
	assert RAM(2260) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(2260))))  severity failure;
	assert RAM(2261) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(2261))))  severity failure;
	assert RAM(2262) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2262))))  severity failure;
	assert RAM(2263) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(2263))))  severity failure;
	assert RAM(2264) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(2264))))  severity failure;
	assert RAM(2265) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2265))))  severity failure;
	assert RAM(2266) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(2266))))  severity failure;
	assert RAM(2267) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(2267))))  severity failure;
	assert RAM(2268) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(2268))))  severity failure;
	assert RAM(2269) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(2269))))  severity failure;
	assert RAM(2270) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(2270))))  severity failure;
	assert RAM(2271) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2271))))  severity failure;
	assert RAM(2272) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(2272))))  severity failure;
	assert RAM(2273) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(2273))))  severity failure;
    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;
end projecttb;
