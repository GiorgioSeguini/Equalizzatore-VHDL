library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
entity project_tb is
end project_tb;
architecture projecttb of project_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;
type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (
			0 => std_logic_vector(to_unsigned(97, 8)),
			1 => std_logic_vector(to_unsigned(120, 8)),
			2 => std_logic_vector(to_unsigned(255, 8)),
			3 => std_logic_vector(to_unsigned(163, 8)),
			4 => std_logic_vector(to_unsigned(111, 8)),
			5 => std_logic_vector(to_unsigned(254, 8)),
			6 => std_logic_vector(to_unsigned(36, 8)),
			7 => std_logic_vector(to_unsigned(60, 8)),
			8 => std_logic_vector(to_unsigned(113, 8)),
			9 => std_logic_vector(to_unsigned(209, 8)),
			10 => std_logic_vector(to_unsigned(194, 8)),
			11 => std_logic_vector(to_unsigned(52, 8)),
			12 => std_logic_vector(to_unsigned(83, 8)),
			13 => std_logic_vector(to_unsigned(215, 8)),
			14 => std_logic_vector(to_unsigned(39, 8)),
			15 => std_logic_vector(to_unsigned(1, 8)),
			16 => std_logic_vector(to_unsigned(8, 8)),
			17 => std_logic_vector(to_unsigned(129, 8)),
			18 => std_logic_vector(to_unsigned(155, 8)),
			19 => std_logic_vector(to_unsigned(173, 8)),
			20 => std_logic_vector(to_unsigned(65, 8)),
			21 => std_logic_vector(to_unsigned(109, 8)),
			22 => std_logic_vector(to_unsigned(183, 8)),
			23 => std_logic_vector(to_unsigned(197, 8)),
			24 => std_logic_vector(to_unsigned(28, 8)),
			25 => std_logic_vector(to_unsigned(188, 8)),
			26 => std_logic_vector(to_unsigned(122, 8)),
			27 => std_logic_vector(to_unsigned(71, 8)),
			28 => std_logic_vector(to_unsigned(114, 8)),
			29 => std_logic_vector(to_unsigned(141, 8)),
			30 => std_logic_vector(to_unsigned(82, 8)),
			31 => std_logic_vector(to_unsigned(85, 8)),
			32 => std_logic_vector(to_unsigned(5, 8)),
			33 => std_logic_vector(to_unsigned(107, 8)),
			34 => std_logic_vector(to_unsigned(74, 8)),
			35 => std_logic_vector(to_unsigned(95, 8)),
			36 => std_logic_vector(to_unsigned(76, 8)),
			37 => std_logic_vector(to_unsigned(80, 8)),
			38 => std_logic_vector(to_unsigned(156, 8)),
			39 => std_logic_vector(to_unsigned(164, 8)),
			40 => std_logic_vector(to_unsigned(181, 8)),
			41 => std_logic_vector(to_unsigned(20, 8)),
			42 => std_logic_vector(to_unsigned(75, 8)),
			43 => std_logic_vector(to_unsigned(113, 8)),
			44 => std_logic_vector(to_unsigned(63, 8)),
			45 => std_logic_vector(to_unsigned(8, 8)),
			46 => std_logic_vector(to_unsigned(129, 8)),
			47 => std_logic_vector(to_unsigned(178, 8)),
			48 => std_logic_vector(to_unsigned(174, 8)),
			49 => std_logic_vector(to_unsigned(91, 8)),
			50 => std_logic_vector(to_unsigned(220, 8)),
			51 => std_logic_vector(to_unsigned(149, 8)),
			52 => std_logic_vector(to_unsigned(255, 8)),
			53 => std_logic_vector(to_unsigned(64, 8)),
			54 => std_logic_vector(to_unsigned(26, 8)),
			55 => std_logic_vector(to_unsigned(12, 8)),
			56 => std_logic_vector(to_unsigned(174, 8)),
			57 => std_logic_vector(to_unsigned(245, 8)),
			58 => std_logic_vector(to_unsigned(133, 8)),
			59 => std_logic_vector(to_unsigned(88, 8)),
			60 => std_logic_vector(to_unsigned(238, 8)),
			61 => std_logic_vector(to_unsigned(53, 8)),
			62 => std_logic_vector(to_unsigned(162, 8)),
			63 => std_logic_vector(to_unsigned(169, 8)),
			64 => std_logic_vector(to_unsigned(9, 8)),
			65 => std_logic_vector(to_unsigned(244, 8)),
			66 => std_logic_vector(to_unsigned(152, 8)),
			67 => std_logic_vector(to_unsigned(210, 8)),
			68 => std_logic_vector(to_unsigned(254, 8)),
			69 => std_logic_vector(to_unsigned(4, 8)),
			70 => std_logic_vector(to_unsigned(86, 8)),
			71 => std_logic_vector(to_unsigned(242, 8)),
			72 => std_logic_vector(to_unsigned(25, 8)),
			73 => std_logic_vector(to_unsigned(230, 8)),
			74 => std_logic_vector(to_unsigned(207, 8)),
			75 => std_logic_vector(to_unsigned(225, 8)),
			76 => std_logic_vector(to_unsigned(80, 8)),
			77 => std_logic_vector(to_unsigned(17, 8)),
			78 => std_logic_vector(to_unsigned(225, 8)),
			79 => std_logic_vector(to_unsigned(116, 8)),
			80 => std_logic_vector(to_unsigned(16, 8)),
			81 => std_logic_vector(to_unsigned(211, 8)),
			82 => std_logic_vector(to_unsigned(254, 8)),
			83 => std_logic_vector(to_unsigned(33, 8)),
			84 => std_logic_vector(to_unsigned(59, 8)),
			85 => std_logic_vector(to_unsigned(79, 8)),
			86 => std_logic_vector(to_unsigned(117, 8)),
			87 => std_logic_vector(to_unsigned(136, 8)),
			88 => std_logic_vector(to_unsigned(2, 8)),
			89 => std_logic_vector(to_unsigned(73, 8)),
			90 => std_logic_vector(to_unsigned(97, 8)),
			91 => std_logic_vector(to_unsigned(186, 8)),
			92 => std_logic_vector(to_unsigned(176, 8)),
			93 => std_logic_vector(to_unsigned(113, 8)),
			94 => std_logic_vector(to_unsigned(207, 8)),
			95 => std_logic_vector(to_unsigned(134, 8)),
			96 => std_logic_vector(to_unsigned(60, 8)),
			97 => std_logic_vector(to_unsigned(196, 8)),
			98 => std_logic_vector(to_unsigned(57, 8)),
			99 => std_logic_vector(to_unsigned(140, 8)),
			100 => std_logic_vector(to_unsigned(239, 8)),
			101 => std_logic_vector(to_unsigned(219, 8)),
			102 => std_logic_vector(to_unsigned(23, 8)),
			103 => std_logic_vector(to_unsigned(221, 8)),
			104 => std_logic_vector(to_unsigned(171, 8)),
			105 => std_logic_vector(to_unsigned(60, 8)),
			106 => std_logic_vector(to_unsigned(249, 8)),
			107 => std_logic_vector(to_unsigned(163, 8)),
			108 => std_logic_vector(to_unsigned(239, 8)),
			109 => std_logic_vector(to_unsigned(205, 8)),
			110 => std_logic_vector(to_unsigned(94, 8)),
			111 => std_logic_vector(to_unsigned(121, 8)),
			112 => std_logic_vector(to_unsigned(70, 8)),
			113 => std_logic_vector(to_unsigned(220, 8)),
			114 => std_logic_vector(to_unsigned(91, 8)),
			115 => std_logic_vector(to_unsigned(232, 8)),
			116 => std_logic_vector(to_unsigned(87, 8)),
			117 => std_logic_vector(to_unsigned(121, 8)),
			118 => std_logic_vector(to_unsigned(155, 8)),
			119 => std_logic_vector(to_unsigned(42, 8)),
			120 => std_logic_vector(to_unsigned(237, 8)),
			121 => std_logic_vector(to_unsigned(92, 8)),
			122 => std_logic_vector(to_unsigned(125, 8)),
			123 => std_logic_vector(to_unsigned(125, 8)),
			124 => std_logic_vector(to_unsigned(243, 8)),
			125 => std_logic_vector(to_unsigned(58, 8)),
			126 => std_logic_vector(to_unsigned(96, 8)),
			127 => std_logic_vector(to_unsigned(160, 8)),
			128 => std_logic_vector(to_unsigned(13, 8)),
			129 => std_logic_vector(to_unsigned(112, 8)),
			130 => std_logic_vector(to_unsigned(237, 8)),
			131 => std_logic_vector(to_unsigned(15, 8)),
			132 => std_logic_vector(to_unsigned(215, 8)),
			133 => std_logic_vector(to_unsigned(206, 8)),
			134 => std_logic_vector(to_unsigned(197, 8)),
			135 => std_logic_vector(to_unsigned(55, 8)),
			136 => std_logic_vector(to_unsigned(144, 8)),
			137 => std_logic_vector(to_unsigned(129, 8)),
			138 => std_logic_vector(to_unsigned(74, 8)),
			139 => std_logic_vector(to_unsigned(103, 8)),
			140 => std_logic_vector(to_unsigned(44, 8)),
			141 => std_logic_vector(to_unsigned(105, 8)),
			142 => std_logic_vector(to_unsigned(33, 8)),
			143 => std_logic_vector(to_unsigned(133, 8)),
			144 => std_logic_vector(to_unsigned(111, 8)),
			145 => std_logic_vector(to_unsigned(230, 8)),
			146 => std_logic_vector(to_unsigned(128, 8)),
			147 => std_logic_vector(to_unsigned(48, 8)),
			148 => std_logic_vector(to_unsigned(22, 8)),
			149 => std_logic_vector(to_unsigned(51, 8)),
			150 => std_logic_vector(to_unsigned(104, 8)),
			151 => std_logic_vector(to_unsigned(129, 8)),
			152 => std_logic_vector(to_unsigned(122, 8)),
			153 => std_logic_vector(to_unsigned(101, 8)),
			154 => std_logic_vector(to_unsigned(147, 8)),
			155 => std_logic_vector(to_unsigned(214, 8)),
			156 => std_logic_vector(to_unsigned(178, 8)),
			157 => std_logic_vector(to_unsigned(130, 8)),
			158 => std_logic_vector(to_unsigned(120, 8)),
			159 => std_logic_vector(to_unsigned(15, 8)),
			160 => std_logic_vector(to_unsigned(59, 8)),
			161 => std_logic_vector(to_unsigned(116, 8)),
			162 => std_logic_vector(to_unsigned(163, 8)),
			163 => std_logic_vector(to_unsigned(243, 8)),
			164 => std_logic_vector(to_unsigned(16, 8)),
			165 => std_logic_vector(to_unsigned(56, 8)),
			166 => std_logic_vector(to_unsigned(84, 8)),
			167 => std_logic_vector(to_unsigned(221, 8)),
			168 => std_logic_vector(to_unsigned(99, 8)),
			169 => std_logic_vector(to_unsigned(196, 8)),
			170 => std_logic_vector(to_unsigned(15, 8)),
			171 => std_logic_vector(to_unsigned(103, 8)),
			172 => std_logic_vector(to_unsigned(168, 8)),
			173 => std_logic_vector(to_unsigned(113, 8)),
			174 => std_logic_vector(to_unsigned(89, 8)),
			175 => std_logic_vector(to_unsigned(40, 8)),
			176 => std_logic_vector(to_unsigned(146, 8)),
			177 => std_logic_vector(to_unsigned(250, 8)),
			178 => std_logic_vector(to_unsigned(12, 8)),
			179 => std_logic_vector(to_unsigned(166, 8)),
			180 => std_logic_vector(to_unsigned(62, 8)),
			181 => std_logic_vector(to_unsigned(250, 8)),
			182 => std_logic_vector(to_unsigned(77, 8)),
			183 => std_logic_vector(to_unsigned(5, 8)),
			184 => std_logic_vector(to_unsigned(80, 8)),
			185 => std_logic_vector(to_unsigned(18, 8)),
			186 => std_logic_vector(to_unsigned(110, 8)),
			187 => std_logic_vector(to_unsigned(60, 8)),
			188 => std_logic_vector(to_unsigned(143, 8)),
			189 => std_logic_vector(to_unsigned(193, 8)),
			190 => std_logic_vector(to_unsigned(117, 8)),
			191 => std_logic_vector(to_unsigned(17, 8)),
			192 => std_logic_vector(to_unsigned(25, 8)),
			193 => std_logic_vector(to_unsigned(170, 8)),
			194 => std_logic_vector(to_unsigned(3, 8)),
			195 => std_logic_vector(to_unsigned(210, 8)),
			196 => std_logic_vector(to_unsigned(8, 8)),
			197 => std_logic_vector(to_unsigned(48, 8)),
			198 => std_logic_vector(to_unsigned(27, 8)),
			199 => std_logic_vector(to_unsigned(12, 8)),
			200 => std_logic_vector(to_unsigned(47, 8)),
			201 => std_logic_vector(to_unsigned(113, 8)),
			202 => std_logic_vector(to_unsigned(95, 8)),
			203 => std_logic_vector(to_unsigned(249, 8)),
			204 => std_logic_vector(to_unsigned(146, 8)),
			205 => std_logic_vector(to_unsigned(78, 8)),
			206 => std_logic_vector(to_unsigned(125, 8)),
			207 => std_logic_vector(to_unsigned(187, 8)),
			208 => std_logic_vector(to_unsigned(91, 8)),
			209 => std_logic_vector(to_unsigned(59, 8)),
			210 => std_logic_vector(to_unsigned(250, 8)),
			211 => std_logic_vector(to_unsigned(225, 8)),
			212 => std_logic_vector(to_unsigned(220, 8)),
			213 => std_logic_vector(to_unsigned(255, 8)),
			214 => std_logic_vector(to_unsigned(24, 8)),
			215 => std_logic_vector(to_unsigned(39, 8)),
			216 => std_logic_vector(to_unsigned(222, 8)),
			217 => std_logic_vector(to_unsigned(168, 8)),
			218 => std_logic_vector(to_unsigned(28, 8)),
			219 => std_logic_vector(to_unsigned(98, 8)),
			220 => std_logic_vector(to_unsigned(146, 8)),
			221 => std_logic_vector(to_unsigned(147, 8)),
			222 => std_logic_vector(to_unsigned(196, 8)),
			223 => std_logic_vector(to_unsigned(222, 8)),
			224 => std_logic_vector(to_unsigned(251, 8)),
			225 => std_logic_vector(to_unsigned(202, 8)),
			226 => std_logic_vector(to_unsigned(141, 8)),
			227 => std_logic_vector(to_unsigned(182, 8)),
			228 => std_logic_vector(to_unsigned(155, 8)),
			229 => std_logic_vector(to_unsigned(216, 8)),
			230 => std_logic_vector(to_unsigned(18, 8)),
			231 => std_logic_vector(to_unsigned(236, 8)),
			232 => std_logic_vector(to_unsigned(208, 8)),
			233 => std_logic_vector(to_unsigned(8, 8)),
			234 => std_logic_vector(to_unsigned(171, 8)),
			235 => std_logic_vector(to_unsigned(173, 8)),
			236 => std_logic_vector(to_unsigned(228, 8)),
			237 => std_logic_vector(to_unsigned(155, 8)),
			238 => std_logic_vector(to_unsigned(92, 8)),
			239 => std_logic_vector(to_unsigned(66, 8)),
			240 => std_logic_vector(to_unsigned(241, 8)),
			241 => std_logic_vector(to_unsigned(59, 8)),
			242 => std_logic_vector(to_unsigned(107, 8)),
			243 => std_logic_vector(to_unsigned(198, 8)),
			244 => std_logic_vector(to_unsigned(244, 8)),
			245 => std_logic_vector(to_unsigned(119, 8)),
			246 => std_logic_vector(to_unsigned(10, 8)),
			247 => std_logic_vector(to_unsigned(94, 8)),
			248 => std_logic_vector(to_unsigned(182, 8)),
			249 => std_logic_vector(to_unsigned(1, 8)),
			250 => std_logic_vector(to_unsigned(71, 8)),
			251 => std_logic_vector(to_unsigned(61, 8)),
			252 => std_logic_vector(to_unsigned(95, 8)),
			253 => std_logic_vector(to_unsigned(73, 8)),
			254 => std_logic_vector(to_unsigned(200, 8)),
			255 => std_logic_vector(to_unsigned(202, 8)),
			256 => std_logic_vector(to_unsigned(131, 8)),
			257 => std_logic_vector(to_unsigned(103, 8)),
			258 => std_logic_vector(to_unsigned(155, 8)),
			259 => std_logic_vector(to_unsigned(185, 8)),
			260 => std_logic_vector(to_unsigned(227, 8)),
			261 => std_logic_vector(to_unsigned(178, 8)),
			262 => std_logic_vector(to_unsigned(251, 8)),
			263 => std_logic_vector(to_unsigned(74, 8)),
			264 => std_logic_vector(to_unsigned(34, 8)),
			265 => std_logic_vector(to_unsigned(124, 8)),
			266 => std_logic_vector(to_unsigned(242, 8)),
			267 => std_logic_vector(to_unsigned(75, 8)),
			268 => std_logic_vector(to_unsigned(1, 8)),
			269 => std_logic_vector(to_unsigned(8, 8)),
			270 => std_logic_vector(to_unsigned(7, 8)),
			271 => std_logic_vector(to_unsigned(75, 8)),
			272 => std_logic_vector(to_unsigned(83, 8)),
			273 => std_logic_vector(to_unsigned(92, 8)),
			274 => std_logic_vector(to_unsigned(40, 8)),
			275 => std_logic_vector(to_unsigned(70, 8)),
			276 => std_logic_vector(to_unsigned(109, 8)),
			277 => std_logic_vector(to_unsigned(224, 8)),
			278 => std_logic_vector(to_unsigned(145, 8)),
			279 => std_logic_vector(to_unsigned(110, 8)),
			280 => std_logic_vector(to_unsigned(227, 8)),
			281 => std_logic_vector(to_unsigned(124, 8)),
			282 => std_logic_vector(to_unsigned(112, 8)),
			283 => std_logic_vector(to_unsigned(167, 8)),
			284 => std_logic_vector(to_unsigned(146, 8)),
			285 => std_logic_vector(to_unsigned(133, 8)),
			286 => std_logic_vector(to_unsigned(80, 8)),
			287 => std_logic_vector(to_unsigned(238, 8)),
			288 => std_logic_vector(to_unsigned(65, 8)),
			289 => std_logic_vector(to_unsigned(197, 8)),
			290 => std_logic_vector(to_unsigned(25, 8)),
			291 => std_logic_vector(to_unsigned(46, 8)),
			292 => std_logic_vector(to_unsigned(208, 8)),
			293 => std_logic_vector(to_unsigned(162, 8)),
			294 => std_logic_vector(to_unsigned(117, 8)),
			295 => std_logic_vector(to_unsigned(14, 8)),
			296 => std_logic_vector(to_unsigned(13, 8)),
			297 => std_logic_vector(to_unsigned(153, 8)),
			298 => std_logic_vector(to_unsigned(188, 8)),
			299 => std_logic_vector(to_unsigned(251, 8)),
			300 => std_logic_vector(to_unsigned(132, 8)),
			301 => std_logic_vector(to_unsigned(78, 8)),
			302 => std_logic_vector(to_unsigned(227, 8)),
			303 => std_logic_vector(to_unsigned(124, 8)),
			304 => std_logic_vector(to_unsigned(169, 8)),
			305 => std_logic_vector(to_unsigned(244, 8)),
			306 => std_logic_vector(to_unsigned(110, 8)),
			307 => std_logic_vector(to_unsigned(160, 8)),
			308 => std_logic_vector(to_unsigned(12, 8)),
			309 => std_logic_vector(to_unsigned(75, 8)),
			310 => std_logic_vector(to_unsigned(32, 8)),
			311 => std_logic_vector(to_unsigned(152, 8)),
			312 => std_logic_vector(to_unsigned(128, 8)),
			313 => std_logic_vector(to_unsigned(73, 8)),
			314 => std_logic_vector(to_unsigned(131, 8)),
			315 => std_logic_vector(to_unsigned(64, 8)),
			316 => std_logic_vector(to_unsigned(98, 8)),
			317 => std_logic_vector(to_unsigned(18, 8)),
			318 => std_logic_vector(to_unsigned(97, 8)),
			319 => std_logic_vector(to_unsigned(18, 8)),
			320 => std_logic_vector(to_unsigned(133, 8)),
			321 => std_logic_vector(to_unsigned(100, 8)),
			322 => std_logic_vector(to_unsigned(67, 8)),
			323 => std_logic_vector(to_unsigned(142, 8)),
			324 => std_logic_vector(to_unsigned(153, 8)),
			325 => std_logic_vector(to_unsigned(253, 8)),
			326 => std_logic_vector(to_unsigned(252, 8)),
			327 => std_logic_vector(to_unsigned(157, 8)),
			328 => std_logic_vector(to_unsigned(212, 8)),
			329 => std_logic_vector(to_unsigned(145, 8)),
			330 => std_logic_vector(to_unsigned(108, 8)),
			331 => std_logic_vector(to_unsigned(97, 8)),
			332 => std_logic_vector(to_unsigned(201, 8)),
			333 => std_logic_vector(to_unsigned(228, 8)),
			334 => std_logic_vector(to_unsigned(61, 8)),
			335 => std_logic_vector(to_unsigned(172, 8)),
			336 => std_logic_vector(to_unsigned(162, 8)),
			337 => std_logic_vector(to_unsigned(39, 8)),
			338 => std_logic_vector(to_unsigned(230, 8)),
			339 => std_logic_vector(to_unsigned(218, 8)),
			340 => std_logic_vector(to_unsigned(236, 8)),
			341 => std_logic_vector(to_unsigned(133, 8)),
			342 => std_logic_vector(to_unsigned(35, 8)),
			343 => std_logic_vector(to_unsigned(148, 8)),
			344 => std_logic_vector(to_unsigned(74, 8)),
			345 => std_logic_vector(to_unsigned(4, 8)),
			346 => std_logic_vector(to_unsigned(172, 8)),
			347 => std_logic_vector(to_unsigned(10, 8)),
			348 => std_logic_vector(to_unsigned(146, 8)),
			349 => std_logic_vector(to_unsigned(26, 8)),
			350 => std_logic_vector(to_unsigned(126, 8)),
			351 => std_logic_vector(to_unsigned(171, 8)),
			352 => std_logic_vector(to_unsigned(6, 8)),
			353 => std_logic_vector(to_unsigned(76, 8)),
			354 => std_logic_vector(to_unsigned(80, 8)),
			355 => std_logic_vector(to_unsigned(167, 8)),
			356 => std_logic_vector(to_unsigned(138, 8)),
			357 => std_logic_vector(to_unsigned(174, 8)),
			358 => std_logic_vector(to_unsigned(34, 8)),
			359 => std_logic_vector(to_unsigned(14, 8)),
			360 => std_logic_vector(to_unsigned(251, 8)),
			361 => std_logic_vector(to_unsigned(218, 8)),
			362 => std_logic_vector(to_unsigned(75, 8)),
			363 => std_logic_vector(to_unsigned(48, 8)),
			364 => std_logic_vector(to_unsigned(41, 8)),
			365 => std_logic_vector(to_unsigned(25, 8)),
			366 => std_logic_vector(to_unsigned(154, 8)),
			367 => std_logic_vector(to_unsigned(51, 8)),
			368 => std_logic_vector(to_unsigned(91, 8)),
			369 => std_logic_vector(to_unsigned(181, 8)),
			370 => std_logic_vector(to_unsigned(72, 8)),
			371 => std_logic_vector(to_unsigned(111, 8)),
			372 => std_logic_vector(to_unsigned(84, 8)),
			373 => std_logic_vector(to_unsigned(192, 8)),
			374 => std_logic_vector(to_unsigned(115, 8)),
			375 => std_logic_vector(to_unsigned(220, 8)),
			376 => std_logic_vector(to_unsigned(73, 8)),
			377 => std_logic_vector(to_unsigned(77, 8)),
			378 => std_logic_vector(to_unsigned(55, 8)),
			379 => std_logic_vector(to_unsigned(111, 8)),
			380 => std_logic_vector(to_unsigned(151, 8)),
			381 => std_logic_vector(to_unsigned(151, 8)),
			382 => std_logic_vector(to_unsigned(235, 8)),
			383 => std_logic_vector(to_unsigned(98, 8)),
			384 => std_logic_vector(to_unsigned(166, 8)),
			385 => std_logic_vector(to_unsigned(180, 8)),
			386 => std_logic_vector(to_unsigned(173, 8)),
			387 => std_logic_vector(to_unsigned(117, 8)),
			388 => std_logic_vector(to_unsigned(89, 8)),
			389 => std_logic_vector(to_unsigned(133, 8)),
			390 => std_logic_vector(to_unsigned(173, 8)),
			391 => std_logic_vector(to_unsigned(175, 8)),
			392 => std_logic_vector(to_unsigned(160, 8)),
			393 => std_logic_vector(to_unsigned(248, 8)),
			394 => std_logic_vector(to_unsigned(26, 8)),
			395 => std_logic_vector(to_unsigned(133, 8)),
			396 => std_logic_vector(to_unsigned(66, 8)),
			397 => std_logic_vector(to_unsigned(255, 8)),
			398 => std_logic_vector(to_unsigned(168, 8)),
			399 => std_logic_vector(to_unsigned(101, 8)),
			400 => std_logic_vector(to_unsigned(86, 8)),
			401 => std_logic_vector(to_unsigned(130, 8)),
			402 => std_logic_vector(to_unsigned(138, 8)),
			403 => std_logic_vector(to_unsigned(103, 8)),
			404 => std_logic_vector(to_unsigned(222, 8)),
			405 => std_logic_vector(to_unsigned(191, 8)),
			406 => std_logic_vector(to_unsigned(197, 8)),
			407 => std_logic_vector(to_unsigned(13, 8)),
			408 => std_logic_vector(to_unsigned(5, 8)),
			409 => std_logic_vector(to_unsigned(81, 8)),
			410 => std_logic_vector(to_unsigned(116, 8)),
			411 => std_logic_vector(to_unsigned(132, 8)),
			412 => std_logic_vector(to_unsigned(53, 8)),
			413 => std_logic_vector(to_unsigned(174, 8)),
			414 => std_logic_vector(to_unsigned(43, 8)),
			415 => std_logic_vector(to_unsigned(175, 8)),
			416 => std_logic_vector(to_unsigned(186, 8)),
			417 => std_logic_vector(to_unsigned(171, 8)),
			418 => std_logic_vector(to_unsigned(231, 8)),
			419 => std_logic_vector(to_unsigned(189, 8)),
			420 => std_logic_vector(to_unsigned(118, 8)),
			421 => std_logic_vector(to_unsigned(182, 8)),
			422 => std_logic_vector(to_unsigned(155, 8)),
			423 => std_logic_vector(to_unsigned(117, 8)),
			424 => std_logic_vector(to_unsigned(238, 8)),
			425 => std_logic_vector(to_unsigned(45, 8)),
			426 => std_logic_vector(to_unsigned(78, 8)),
			427 => std_logic_vector(to_unsigned(74, 8)),
			428 => std_logic_vector(to_unsigned(77, 8)),
			429 => std_logic_vector(to_unsigned(220, 8)),
			430 => std_logic_vector(to_unsigned(145, 8)),
			431 => std_logic_vector(to_unsigned(189, 8)),
			432 => std_logic_vector(to_unsigned(39, 8)),
			433 => std_logic_vector(to_unsigned(152, 8)),
			434 => std_logic_vector(to_unsigned(136, 8)),
			435 => std_logic_vector(to_unsigned(171, 8)),
			436 => std_logic_vector(to_unsigned(181, 8)),
			437 => std_logic_vector(to_unsigned(136, 8)),
			438 => std_logic_vector(to_unsigned(234, 8)),
			439 => std_logic_vector(to_unsigned(196, 8)),
			440 => std_logic_vector(to_unsigned(196, 8)),
			441 => std_logic_vector(to_unsigned(57, 8)),
			442 => std_logic_vector(to_unsigned(217, 8)),
			443 => std_logic_vector(to_unsigned(219, 8)),
			444 => std_logic_vector(to_unsigned(13, 8)),
			445 => std_logic_vector(to_unsigned(126, 8)),
			446 => std_logic_vector(to_unsigned(2, 8)),
			447 => std_logic_vector(to_unsigned(81, 8)),
			448 => std_logic_vector(to_unsigned(4, 8)),
			449 => std_logic_vector(to_unsigned(251, 8)),
			450 => std_logic_vector(to_unsigned(121, 8)),
			451 => std_logic_vector(to_unsigned(140, 8)),
			452 => std_logic_vector(to_unsigned(178, 8)),
			453 => std_logic_vector(to_unsigned(235, 8)),
			454 => std_logic_vector(to_unsigned(246, 8)),
			455 => std_logic_vector(to_unsigned(16, 8)),
			456 => std_logic_vector(to_unsigned(51, 8)),
			457 => std_logic_vector(to_unsigned(194, 8)),
			458 => std_logic_vector(to_unsigned(93, 8)),
			459 => std_logic_vector(to_unsigned(226, 8)),
			460 => std_logic_vector(to_unsigned(40, 8)),
			461 => std_logic_vector(to_unsigned(23, 8)),
			462 => std_logic_vector(to_unsigned(64, 8)),
			463 => std_logic_vector(to_unsigned(164, 8)),
			464 => std_logic_vector(to_unsigned(186, 8)),
			465 => std_logic_vector(to_unsigned(126, 8)),
			466 => std_logic_vector(to_unsigned(235, 8)),
			467 => std_logic_vector(to_unsigned(202, 8)),
			468 => std_logic_vector(to_unsigned(31, 8)),
			469 => std_logic_vector(to_unsigned(147, 8)),
			470 => std_logic_vector(to_unsigned(81, 8)),
			471 => std_logic_vector(to_unsigned(121, 8)),
			472 => std_logic_vector(to_unsigned(238, 8)),
			473 => std_logic_vector(to_unsigned(7, 8)),
			474 => std_logic_vector(to_unsigned(20, 8)),
			475 => std_logic_vector(to_unsigned(130, 8)),
			476 => std_logic_vector(to_unsigned(9, 8)),
			477 => std_logic_vector(to_unsigned(34, 8)),
			478 => std_logic_vector(to_unsigned(140, 8)),
			479 => std_logic_vector(to_unsigned(63, 8)),
			480 => std_logic_vector(to_unsigned(10, 8)),
			481 => std_logic_vector(to_unsigned(36, 8)),
			482 => std_logic_vector(to_unsigned(208, 8)),
			483 => std_logic_vector(to_unsigned(105, 8)),
			484 => std_logic_vector(to_unsigned(174, 8)),
			485 => std_logic_vector(to_unsigned(105, 8)),
			486 => std_logic_vector(to_unsigned(224, 8)),
			487 => std_logic_vector(to_unsigned(205, 8)),
			488 => std_logic_vector(to_unsigned(7, 8)),
			489 => std_logic_vector(to_unsigned(12, 8)),
			490 => std_logic_vector(to_unsigned(85, 8)),
			491 => std_logic_vector(to_unsigned(100, 8)),
			492 => std_logic_vector(to_unsigned(223, 8)),
			493 => std_logic_vector(to_unsigned(161, 8)),
			494 => std_logic_vector(to_unsigned(176, 8)),
			495 => std_logic_vector(to_unsigned(230, 8)),
			496 => std_logic_vector(to_unsigned(165, 8)),
			497 => std_logic_vector(to_unsigned(99, 8)),
			498 => std_logic_vector(to_unsigned(216, 8)),
			499 => std_logic_vector(to_unsigned(142, 8)),
			500 => std_logic_vector(to_unsigned(122, 8)),
			501 => std_logic_vector(to_unsigned(35, 8)),
			502 => std_logic_vector(to_unsigned(194, 8)),
			503 => std_logic_vector(to_unsigned(112, 8)),
			504 => std_logic_vector(to_unsigned(190, 8)),
			505 => std_logic_vector(to_unsigned(243, 8)),
			506 => std_logic_vector(to_unsigned(41, 8)),
			507 => std_logic_vector(to_unsigned(51, 8)),
			508 => std_logic_vector(to_unsigned(37, 8)),
			509 => std_logic_vector(to_unsigned(192, 8)),
			510 => std_logic_vector(to_unsigned(197, 8)),
			511 => std_logic_vector(to_unsigned(82, 8)),
			512 => std_logic_vector(to_unsigned(91, 8)),
			513 => std_logic_vector(to_unsigned(120, 8)),
			514 => std_logic_vector(to_unsigned(143, 8)),
			515 => std_logic_vector(to_unsigned(99, 8)),
			516 => std_logic_vector(to_unsigned(239, 8)),
			517 => std_logic_vector(to_unsigned(139, 8)),
			518 => std_logic_vector(to_unsigned(205, 8)),
			519 => std_logic_vector(to_unsigned(69, 8)),
			520 => std_logic_vector(to_unsigned(198, 8)),
			521 => std_logic_vector(to_unsigned(36, 8)),
			522 => std_logic_vector(to_unsigned(192, 8)),
			523 => std_logic_vector(to_unsigned(252, 8)),
			524 => std_logic_vector(to_unsigned(6, 8)),
			525 => std_logic_vector(to_unsigned(2, 8)),
			526 => std_logic_vector(to_unsigned(206, 8)),
			527 => std_logic_vector(to_unsigned(253, 8)),
			528 => std_logic_vector(to_unsigned(85, 8)),
			529 => std_logic_vector(to_unsigned(46, 8)),
			530 => std_logic_vector(to_unsigned(254, 8)),
			531 => std_logic_vector(to_unsigned(202, 8)),
			532 => std_logic_vector(to_unsigned(120, 8)),
			533 => std_logic_vector(to_unsigned(248, 8)),
			534 => std_logic_vector(to_unsigned(84, 8)),
			535 => std_logic_vector(to_unsigned(146, 8)),
			536 => std_logic_vector(to_unsigned(175, 8)),
			537 => std_logic_vector(to_unsigned(168, 8)),
			538 => std_logic_vector(to_unsigned(225, 8)),
			539 => std_logic_vector(to_unsigned(58, 8)),
			540 => std_logic_vector(to_unsigned(197, 8)),
			541 => std_logic_vector(to_unsigned(121, 8)),
			542 => std_logic_vector(to_unsigned(109, 8)),
			543 => std_logic_vector(to_unsigned(177, 8)),
			544 => std_logic_vector(to_unsigned(163, 8)),
			545 => std_logic_vector(to_unsigned(153, 8)),
			546 => std_logic_vector(to_unsigned(188, 8)),
			547 => std_logic_vector(to_unsigned(7, 8)),
			548 => std_logic_vector(to_unsigned(212, 8)),
			549 => std_logic_vector(to_unsigned(168, 8)),
			550 => std_logic_vector(to_unsigned(10, 8)),
			551 => std_logic_vector(to_unsigned(199, 8)),
			552 => std_logic_vector(to_unsigned(48, 8)),
			553 => std_logic_vector(to_unsigned(30, 8)),
			554 => std_logic_vector(to_unsigned(215, 8)),
			555 => std_logic_vector(to_unsigned(62, 8)),
			556 => std_logic_vector(to_unsigned(222, 8)),
			557 => std_logic_vector(to_unsigned(92, 8)),
			558 => std_logic_vector(to_unsigned(7, 8)),
			559 => std_logic_vector(to_unsigned(41, 8)),
			560 => std_logic_vector(to_unsigned(47, 8)),
			561 => std_logic_vector(to_unsigned(178, 8)),
			562 => std_logic_vector(to_unsigned(213, 8)),
			563 => std_logic_vector(to_unsigned(8, 8)),
			564 => std_logic_vector(to_unsigned(210, 8)),
			565 => std_logic_vector(to_unsigned(62, 8)),
			566 => std_logic_vector(to_unsigned(87, 8)),
			567 => std_logic_vector(to_unsigned(233, 8)),
			568 => std_logic_vector(to_unsigned(247, 8)),
			569 => std_logic_vector(to_unsigned(37, 8)),
			570 => std_logic_vector(to_unsigned(217, 8)),
			571 => std_logic_vector(to_unsigned(19, 8)),
			572 => std_logic_vector(to_unsigned(195, 8)),
			573 => std_logic_vector(to_unsigned(19, 8)),
			574 => std_logic_vector(to_unsigned(42, 8)),
			575 => std_logic_vector(to_unsigned(50, 8)),
			576 => std_logic_vector(to_unsigned(219, 8)),
			577 => std_logic_vector(to_unsigned(202, 8)),
			578 => std_logic_vector(to_unsigned(36, 8)),
			579 => std_logic_vector(to_unsigned(129, 8)),
			580 => std_logic_vector(to_unsigned(38, 8)),
			581 => std_logic_vector(to_unsigned(241, 8)),
			582 => std_logic_vector(to_unsigned(88, 8)),
			583 => std_logic_vector(to_unsigned(195, 8)),
			584 => std_logic_vector(to_unsigned(38, 8)),
			585 => std_logic_vector(to_unsigned(99, 8)),
			586 => std_logic_vector(to_unsigned(122, 8)),
			587 => std_logic_vector(to_unsigned(203, 8)),
			588 => std_logic_vector(to_unsigned(158, 8)),
			589 => std_logic_vector(to_unsigned(7, 8)),
			590 => std_logic_vector(to_unsigned(223, 8)),
			591 => std_logic_vector(to_unsigned(31, 8)),
			592 => std_logic_vector(to_unsigned(183, 8)),
			593 => std_logic_vector(to_unsigned(203, 8)),
			594 => std_logic_vector(to_unsigned(244, 8)),
			595 => std_logic_vector(to_unsigned(39, 8)),
			596 => std_logic_vector(to_unsigned(191, 8)),
			597 => std_logic_vector(to_unsigned(78, 8)),
			598 => std_logic_vector(to_unsigned(202, 8)),
			599 => std_logic_vector(to_unsigned(119, 8)),
			600 => std_logic_vector(to_unsigned(118, 8)),
			601 => std_logic_vector(to_unsigned(202, 8)),
			602 => std_logic_vector(to_unsigned(185, 8)),
			603 => std_logic_vector(to_unsigned(108, 8)),
			604 => std_logic_vector(to_unsigned(81, 8)),
			605 => std_logic_vector(to_unsigned(126, 8)),
			606 => std_logic_vector(to_unsigned(34, 8)),
			607 => std_logic_vector(to_unsigned(48, 8)),
			608 => std_logic_vector(to_unsigned(32, 8)),
			609 => std_logic_vector(to_unsigned(19, 8)),
			610 => std_logic_vector(to_unsigned(231, 8)),
			611 => std_logic_vector(to_unsigned(90, 8)),
			612 => std_logic_vector(to_unsigned(149, 8)),
			613 => std_logic_vector(to_unsigned(135, 8)),
			614 => std_logic_vector(to_unsigned(78, 8)),
			615 => std_logic_vector(to_unsigned(118, 8)),
			616 => std_logic_vector(to_unsigned(179, 8)),
			617 => std_logic_vector(to_unsigned(212, 8)),
			618 => std_logic_vector(to_unsigned(74, 8)),
			619 => std_logic_vector(to_unsigned(197, 8)),
			620 => std_logic_vector(to_unsigned(218, 8)),
			621 => std_logic_vector(to_unsigned(113, 8)),
			622 => std_logic_vector(to_unsigned(63, 8)),
			623 => std_logic_vector(to_unsigned(46, 8)),
			624 => std_logic_vector(to_unsigned(68, 8)),
			625 => std_logic_vector(to_unsigned(198, 8)),
			626 => std_logic_vector(to_unsigned(7, 8)),
			627 => std_logic_vector(to_unsigned(52, 8)),
			628 => std_logic_vector(to_unsigned(124, 8)),
			629 => std_logic_vector(to_unsigned(143, 8)),
			630 => std_logic_vector(to_unsigned(241, 8)),
			631 => std_logic_vector(to_unsigned(96, 8)),
			632 => std_logic_vector(to_unsigned(221, 8)),
			633 => std_logic_vector(to_unsigned(102, 8)),
			634 => std_logic_vector(to_unsigned(94, 8)),
			635 => std_logic_vector(to_unsigned(145, 8)),
			636 => std_logic_vector(to_unsigned(184, 8)),
			637 => std_logic_vector(to_unsigned(70, 8)),
			638 => std_logic_vector(to_unsigned(61, 8)),
			639 => std_logic_vector(to_unsigned(213, 8)),
			640 => std_logic_vector(to_unsigned(209, 8)),
			641 => std_logic_vector(to_unsigned(231, 8)),
			642 => std_logic_vector(to_unsigned(8, 8)),
			643 => std_logic_vector(to_unsigned(171, 8)),
			644 => std_logic_vector(to_unsigned(121, 8)),
			645 => std_logic_vector(to_unsigned(180, 8)),
			646 => std_logic_vector(to_unsigned(96, 8)),
			647 => std_logic_vector(to_unsigned(211, 8)),
			648 => std_logic_vector(to_unsigned(7, 8)),
			649 => std_logic_vector(to_unsigned(191, 8)),
			650 => std_logic_vector(to_unsigned(166, 8)),
			651 => std_logic_vector(to_unsigned(19, 8)),
			652 => std_logic_vector(to_unsigned(15, 8)),
			653 => std_logic_vector(to_unsigned(179, 8)),
			654 => std_logic_vector(to_unsigned(250, 8)),
			655 => std_logic_vector(to_unsigned(45, 8)),
			656 => std_logic_vector(to_unsigned(228, 8)),
			657 => std_logic_vector(to_unsigned(189, 8)),
			658 => std_logic_vector(to_unsigned(205, 8)),
			659 => std_logic_vector(to_unsigned(214, 8)),
			660 => std_logic_vector(to_unsigned(210, 8)),
			661 => std_logic_vector(to_unsigned(28, 8)),
			662 => std_logic_vector(to_unsigned(182, 8)),
			663 => std_logic_vector(to_unsigned(81, 8)),
			664 => std_logic_vector(to_unsigned(220, 8)),
			665 => std_logic_vector(to_unsigned(253, 8)),
			666 => std_logic_vector(to_unsigned(152, 8)),
			667 => std_logic_vector(to_unsigned(181, 8)),
			668 => std_logic_vector(to_unsigned(148, 8)),
			669 => std_logic_vector(to_unsigned(163, 8)),
			670 => std_logic_vector(to_unsigned(163, 8)),
			671 => std_logic_vector(to_unsigned(124, 8)),
			672 => std_logic_vector(to_unsigned(117, 8)),
			673 => std_logic_vector(to_unsigned(129, 8)),
			674 => std_logic_vector(to_unsigned(189, 8)),
			675 => std_logic_vector(to_unsigned(23, 8)),
			676 => std_logic_vector(to_unsigned(176, 8)),
			677 => std_logic_vector(to_unsigned(10, 8)),
			678 => std_logic_vector(to_unsigned(67, 8)),
			679 => std_logic_vector(to_unsigned(5, 8)),
			680 => std_logic_vector(to_unsigned(156, 8)),
			681 => std_logic_vector(to_unsigned(213, 8)),
			682 => std_logic_vector(to_unsigned(82, 8)),
			683 => std_logic_vector(to_unsigned(128, 8)),
			684 => std_logic_vector(to_unsigned(115, 8)),
			685 => std_logic_vector(to_unsigned(8, 8)),
			686 => std_logic_vector(to_unsigned(110, 8)),
			687 => std_logic_vector(to_unsigned(109, 8)),
			688 => std_logic_vector(to_unsigned(243, 8)),
			689 => std_logic_vector(to_unsigned(125, 8)),
			690 => std_logic_vector(to_unsigned(15, 8)),
			691 => std_logic_vector(to_unsigned(73, 8)),
			692 => std_logic_vector(to_unsigned(23, 8)),
			693 => std_logic_vector(to_unsigned(246, 8)),
			694 => std_logic_vector(to_unsigned(206, 8)),
			695 => std_logic_vector(to_unsigned(133, 8)),
			696 => std_logic_vector(to_unsigned(66, 8)),
			697 => std_logic_vector(to_unsigned(201, 8)),
			698 => std_logic_vector(to_unsigned(226, 8)),
			699 => std_logic_vector(to_unsigned(146, 8)),
			700 => std_logic_vector(to_unsigned(93, 8)),
			701 => std_logic_vector(to_unsigned(231, 8)),
			702 => std_logic_vector(to_unsigned(173, 8)),
			703 => std_logic_vector(to_unsigned(206, 8)),
			704 => std_logic_vector(to_unsigned(210, 8)),
			705 => std_logic_vector(to_unsigned(181, 8)),
			706 => std_logic_vector(to_unsigned(44, 8)),
			707 => std_logic_vector(to_unsigned(146, 8)),
			708 => std_logic_vector(to_unsigned(102, 8)),
			709 => std_logic_vector(to_unsigned(157, 8)),
			710 => std_logic_vector(to_unsigned(156, 8)),
			711 => std_logic_vector(to_unsigned(52, 8)),
			712 => std_logic_vector(to_unsigned(79, 8)),
			713 => std_logic_vector(to_unsigned(230, 8)),
			714 => std_logic_vector(to_unsigned(202, 8)),
			715 => std_logic_vector(to_unsigned(90, 8)),
			716 => std_logic_vector(to_unsigned(252, 8)),
			717 => std_logic_vector(to_unsigned(127, 8)),
			718 => std_logic_vector(to_unsigned(82, 8)),
			719 => std_logic_vector(to_unsigned(254, 8)),
			720 => std_logic_vector(to_unsigned(139, 8)),
			721 => std_logic_vector(to_unsigned(84, 8)),
			722 => std_logic_vector(to_unsigned(203, 8)),
			723 => std_logic_vector(to_unsigned(249, 8)),
			724 => std_logic_vector(to_unsigned(201, 8)),
			725 => std_logic_vector(to_unsigned(108, 8)),
			726 => std_logic_vector(to_unsigned(10, 8)),
			727 => std_logic_vector(to_unsigned(124, 8)),
			728 => std_logic_vector(to_unsigned(190, 8)),
			729 => std_logic_vector(to_unsigned(138, 8)),
			730 => std_logic_vector(to_unsigned(178, 8)),
			731 => std_logic_vector(to_unsigned(81, 8)),
			732 => std_logic_vector(to_unsigned(235, 8)),
			733 => std_logic_vector(to_unsigned(161, 8)),
			734 => std_logic_vector(to_unsigned(13, 8)),
			735 => std_logic_vector(to_unsigned(89, 8)),
			736 => std_logic_vector(to_unsigned(241, 8)),
			737 => std_logic_vector(to_unsigned(159, 8)),
			738 => std_logic_vector(to_unsigned(177, 8)),
			739 => std_logic_vector(to_unsigned(253, 8)),
			740 => std_logic_vector(to_unsigned(1, 8)),
			741 => std_logic_vector(to_unsigned(93, 8)),
			742 => std_logic_vector(to_unsigned(131, 8)),
			743 => std_logic_vector(to_unsigned(233, 8)),
			744 => std_logic_vector(to_unsigned(121, 8)),
			745 => std_logic_vector(to_unsigned(247, 8)),
			746 => std_logic_vector(to_unsigned(87, 8)),
			747 => std_logic_vector(to_unsigned(197, 8)),
			748 => std_logic_vector(to_unsigned(137, 8)),
			749 => std_logic_vector(to_unsigned(38, 8)),
			750 => std_logic_vector(to_unsigned(157, 8)),
			751 => std_logic_vector(to_unsigned(67, 8)),
			752 => std_logic_vector(to_unsigned(104, 8)),
			753 => std_logic_vector(to_unsigned(118, 8)),
			754 => std_logic_vector(to_unsigned(190, 8)),
			755 => std_logic_vector(to_unsigned(101, 8)),
			756 => std_logic_vector(to_unsigned(70, 8)),
			757 => std_logic_vector(to_unsigned(38, 8)),
			758 => std_logic_vector(to_unsigned(15, 8)),
			759 => std_logic_vector(to_unsigned(179, 8)),
			760 => std_logic_vector(to_unsigned(1, 8)),
			761 => std_logic_vector(to_unsigned(131, 8)),
			762 => std_logic_vector(to_unsigned(152, 8)),
			763 => std_logic_vector(to_unsigned(223, 8)),
			764 => std_logic_vector(to_unsigned(168, 8)),
			765 => std_logic_vector(to_unsigned(209, 8)),
			766 => std_logic_vector(to_unsigned(212, 8)),
			767 => std_logic_vector(to_unsigned(77, 8)),
			768 => std_logic_vector(to_unsigned(217, 8)),
			769 => std_logic_vector(to_unsigned(71, 8)),
			770 => std_logic_vector(to_unsigned(146, 8)),
			771 => std_logic_vector(to_unsigned(67, 8)),
			772 => std_logic_vector(to_unsigned(186, 8)),
			773 => std_logic_vector(to_unsigned(121, 8)),
			774 => std_logic_vector(to_unsigned(87, 8)),
			775 => std_logic_vector(to_unsigned(213, 8)),
			776 => std_logic_vector(to_unsigned(254, 8)),
			777 => std_logic_vector(to_unsigned(235, 8)),
			778 => std_logic_vector(to_unsigned(165, 8)),
			779 => std_logic_vector(to_unsigned(226, 8)),
			780 => std_logic_vector(to_unsigned(226, 8)),
			781 => std_logic_vector(to_unsigned(150, 8)),
			782 => std_logic_vector(to_unsigned(128, 8)),
			783 => std_logic_vector(to_unsigned(108, 8)),
			784 => std_logic_vector(to_unsigned(24, 8)),
			785 => std_logic_vector(to_unsigned(28, 8)),
			786 => std_logic_vector(to_unsigned(250, 8)),
			787 => std_logic_vector(to_unsigned(234, 8)),
			788 => std_logic_vector(to_unsigned(84, 8)),
			789 => std_logic_vector(to_unsigned(82, 8)),
			790 => std_logic_vector(to_unsigned(199, 8)),
			791 => std_logic_vector(to_unsigned(13, 8)),
			792 => std_logic_vector(to_unsigned(188, 8)),
			793 => std_logic_vector(to_unsigned(237, 8)),
			794 => std_logic_vector(to_unsigned(67, 8)),
			795 => std_logic_vector(to_unsigned(5, 8)),
			796 => std_logic_vector(to_unsigned(122, 8)),
			797 => std_logic_vector(to_unsigned(65, 8)),
			798 => std_logic_vector(to_unsigned(6, 8)),
			799 => std_logic_vector(to_unsigned(33, 8)),
			800 => std_logic_vector(to_unsigned(90, 8)),
			801 => std_logic_vector(to_unsigned(81, 8)),
			802 => std_logic_vector(to_unsigned(61, 8)),
			803 => std_logic_vector(to_unsigned(152, 8)),
			804 => std_logic_vector(to_unsigned(40, 8)),
			805 => std_logic_vector(to_unsigned(149, 8)),
			806 => std_logic_vector(to_unsigned(26, 8)),
			807 => std_logic_vector(to_unsigned(241, 8)),
			808 => std_logic_vector(to_unsigned(108, 8)),
			809 => std_logic_vector(to_unsigned(186, 8)),
			810 => std_logic_vector(to_unsigned(92, 8)),
			811 => std_logic_vector(to_unsigned(163, 8)),
			812 => std_logic_vector(to_unsigned(253, 8)),
			813 => std_logic_vector(to_unsigned(245, 8)),
			814 => std_logic_vector(to_unsigned(7, 8)),
			815 => std_logic_vector(to_unsigned(79, 8)),
			816 => std_logic_vector(to_unsigned(130, 8)),
			817 => std_logic_vector(to_unsigned(153, 8)),
			818 => std_logic_vector(to_unsigned(29, 8)),
			819 => std_logic_vector(to_unsigned(128, 8)),
			820 => std_logic_vector(to_unsigned(99, 8)),
			821 => std_logic_vector(to_unsigned(157, 8)),
			822 => std_logic_vector(to_unsigned(112, 8)),
			823 => std_logic_vector(to_unsigned(86, 8)),
			824 => std_logic_vector(to_unsigned(86, 8)),
			825 => std_logic_vector(to_unsigned(69, 8)),
			826 => std_logic_vector(to_unsigned(96, 8)),
			827 => std_logic_vector(to_unsigned(108, 8)),
			828 => std_logic_vector(to_unsigned(66, 8)),
			829 => std_logic_vector(to_unsigned(147, 8)),
			830 => std_logic_vector(to_unsigned(94, 8)),
			831 => std_logic_vector(to_unsigned(238, 8)),
			832 => std_logic_vector(to_unsigned(6, 8)),
			833 => std_logic_vector(to_unsigned(237, 8)),
			834 => std_logic_vector(to_unsigned(237, 8)),
			835 => std_logic_vector(to_unsigned(167, 8)),
			836 => std_logic_vector(to_unsigned(81, 8)),
			837 => std_logic_vector(to_unsigned(47, 8)),
			838 => std_logic_vector(to_unsigned(0, 8)),
			839 => std_logic_vector(to_unsigned(172, 8)),
			840 => std_logic_vector(to_unsigned(74, 8)),
			841 => std_logic_vector(to_unsigned(189, 8)),
			842 => std_logic_vector(to_unsigned(199, 8)),
			843 => std_logic_vector(to_unsigned(67, 8)),
			844 => std_logic_vector(to_unsigned(14, 8)),
			845 => std_logic_vector(to_unsigned(103, 8)),
			846 => std_logic_vector(to_unsigned(76, 8)),
			847 => std_logic_vector(to_unsigned(143, 8)),
			848 => std_logic_vector(to_unsigned(103, 8)),
			849 => std_logic_vector(to_unsigned(178, 8)),
			850 => std_logic_vector(to_unsigned(39, 8)),
			851 => std_logic_vector(to_unsigned(116, 8)),
			852 => std_logic_vector(to_unsigned(138, 8)),
			853 => std_logic_vector(to_unsigned(83, 8)),
			854 => std_logic_vector(to_unsigned(57, 8)),
			855 => std_logic_vector(to_unsigned(105, 8)),
			856 => std_logic_vector(to_unsigned(240, 8)),
			857 => std_logic_vector(to_unsigned(128, 8)),
			858 => std_logic_vector(to_unsigned(11, 8)),
			859 => std_logic_vector(to_unsigned(194, 8)),
			860 => std_logic_vector(to_unsigned(209, 8)),
			861 => std_logic_vector(to_unsigned(238, 8)),
			862 => std_logic_vector(to_unsigned(209, 8)),
			863 => std_logic_vector(to_unsigned(41, 8)),
			864 => std_logic_vector(to_unsigned(93, 8)),
			865 => std_logic_vector(to_unsigned(194, 8)),
			866 => std_logic_vector(to_unsigned(203, 8)),
			867 => std_logic_vector(to_unsigned(92, 8)),
			868 => std_logic_vector(to_unsigned(70, 8)),
			869 => std_logic_vector(to_unsigned(35, 8)),
			870 => std_logic_vector(to_unsigned(122, 8)),
			871 => std_logic_vector(to_unsigned(214, 8)),
			872 => std_logic_vector(to_unsigned(99, 8)),
			873 => std_logic_vector(to_unsigned(139, 8)),
			874 => std_logic_vector(to_unsigned(191, 8)),
			875 => std_logic_vector(to_unsigned(9, 8)),
			876 => std_logic_vector(to_unsigned(12, 8)),
			877 => std_logic_vector(to_unsigned(240, 8)),
			878 => std_logic_vector(to_unsigned(41, 8)),
			879 => std_logic_vector(to_unsigned(54, 8)),
			880 => std_logic_vector(to_unsigned(19, 8)),
			881 => std_logic_vector(to_unsigned(4, 8)),
			882 => std_logic_vector(to_unsigned(51, 8)),
			883 => std_logic_vector(to_unsigned(82, 8)),
			884 => std_logic_vector(to_unsigned(37, 8)),
			885 => std_logic_vector(to_unsigned(141, 8)),
			886 => std_logic_vector(to_unsigned(29, 8)),
			887 => std_logic_vector(to_unsigned(92, 8)),
			888 => std_logic_vector(to_unsigned(247, 8)),
			889 => std_logic_vector(to_unsigned(56, 8)),
			890 => std_logic_vector(to_unsigned(81, 8)),
			891 => std_logic_vector(to_unsigned(206, 8)),
			892 => std_logic_vector(to_unsigned(22, 8)),
			893 => std_logic_vector(to_unsigned(105, 8)),
			894 => std_logic_vector(to_unsigned(68, 8)),
			895 => std_logic_vector(to_unsigned(215, 8)),
			896 => std_logic_vector(to_unsigned(142, 8)),
			897 => std_logic_vector(to_unsigned(155, 8)),
			898 => std_logic_vector(to_unsigned(160, 8)),
			899 => std_logic_vector(to_unsigned(49, 8)),
			900 => std_logic_vector(to_unsigned(100, 8)),
			901 => std_logic_vector(to_unsigned(42, 8)),
			902 => std_logic_vector(to_unsigned(157, 8)),
			903 => std_logic_vector(to_unsigned(65, 8)),
			904 => std_logic_vector(to_unsigned(96, 8)),
			905 => std_logic_vector(to_unsigned(119, 8)),
			906 => std_logic_vector(to_unsigned(214, 8)),
			907 => std_logic_vector(to_unsigned(13, 8)),
			908 => std_logic_vector(to_unsigned(31, 8)),
			909 => std_logic_vector(to_unsigned(146, 8)),
			910 => std_logic_vector(to_unsigned(122, 8)),
			911 => std_logic_vector(to_unsigned(104, 8)),
			912 => std_logic_vector(to_unsigned(187, 8)),
			913 => std_logic_vector(to_unsigned(29, 8)),
			914 => std_logic_vector(to_unsigned(112, 8)),
			915 => std_logic_vector(to_unsigned(225, 8)),
			916 => std_logic_vector(to_unsigned(196, 8)),
			917 => std_logic_vector(to_unsigned(30, 8)),
			918 => std_logic_vector(to_unsigned(161, 8)),
			919 => std_logic_vector(to_unsigned(24, 8)),
			920 => std_logic_vector(to_unsigned(110, 8)),
			921 => std_logic_vector(to_unsigned(78, 8)),
			922 => std_logic_vector(to_unsigned(201, 8)),
			923 => std_logic_vector(to_unsigned(215, 8)),
			924 => std_logic_vector(to_unsigned(24, 8)),
			925 => std_logic_vector(to_unsigned(217, 8)),
			926 => std_logic_vector(to_unsigned(250, 8)),
			927 => std_logic_vector(to_unsigned(151, 8)),
			928 => std_logic_vector(to_unsigned(23, 8)),
			929 => std_logic_vector(to_unsigned(208, 8)),
			930 => std_logic_vector(to_unsigned(30, 8)),
			931 => std_logic_vector(to_unsigned(234, 8)),
			932 => std_logic_vector(to_unsigned(123, 8)),
			933 => std_logic_vector(to_unsigned(89, 8)),
			934 => std_logic_vector(to_unsigned(56, 8)),
			935 => std_logic_vector(to_unsigned(18, 8)),
			936 => std_logic_vector(to_unsigned(244, 8)),
			937 => std_logic_vector(to_unsigned(146, 8)),
			938 => std_logic_vector(to_unsigned(152, 8)),
			939 => std_logic_vector(to_unsigned(37, 8)),
			940 => std_logic_vector(to_unsigned(48, 8)),
			941 => std_logic_vector(to_unsigned(106, 8)),
			942 => std_logic_vector(to_unsigned(5, 8)),
			943 => std_logic_vector(to_unsigned(210, 8)),
			944 => std_logic_vector(to_unsigned(128, 8)),
			945 => std_logic_vector(to_unsigned(151, 8)),
			946 => std_logic_vector(to_unsigned(251, 8)),
			947 => std_logic_vector(to_unsigned(89, 8)),
			948 => std_logic_vector(to_unsigned(6, 8)),
			949 => std_logic_vector(to_unsigned(137, 8)),
			950 => std_logic_vector(to_unsigned(163, 8)),
			951 => std_logic_vector(to_unsigned(187, 8)),
			952 => std_logic_vector(to_unsigned(121, 8)),
			953 => std_logic_vector(to_unsigned(232, 8)),
			954 => std_logic_vector(to_unsigned(65, 8)),
			955 => std_logic_vector(to_unsigned(117, 8)),
			956 => std_logic_vector(to_unsigned(186, 8)),
			957 => std_logic_vector(to_unsigned(250, 8)),
			958 => std_logic_vector(to_unsigned(54, 8)),
			959 => std_logic_vector(to_unsigned(28, 8)),
			960 => std_logic_vector(to_unsigned(219, 8)),
			961 => std_logic_vector(to_unsigned(99, 8)),
			962 => std_logic_vector(to_unsigned(65, 8)),
			963 => std_logic_vector(to_unsigned(36, 8)),
			964 => std_logic_vector(to_unsigned(129, 8)),
			965 => std_logic_vector(to_unsigned(117, 8)),
			966 => std_logic_vector(to_unsigned(127, 8)),
			967 => std_logic_vector(to_unsigned(234, 8)),
			968 => std_logic_vector(to_unsigned(124, 8)),
			969 => std_logic_vector(to_unsigned(49, 8)),
			970 => std_logic_vector(to_unsigned(3, 8)),
			971 => std_logic_vector(to_unsigned(176, 8)),
			972 => std_logic_vector(to_unsigned(230, 8)),
			973 => std_logic_vector(to_unsigned(109, 8)),
			974 => std_logic_vector(to_unsigned(57, 8)),
			975 => std_logic_vector(to_unsigned(231, 8)),
			976 => std_logic_vector(to_unsigned(19, 8)),
			977 => std_logic_vector(to_unsigned(240, 8)),
			978 => std_logic_vector(to_unsigned(116, 8)),
			979 => std_logic_vector(to_unsigned(3, 8)),
			980 => std_logic_vector(to_unsigned(8, 8)),
			981 => std_logic_vector(to_unsigned(30, 8)),
			982 => std_logic_vector(to_unsigned(121, 8)),
			983 => std_logic_vector(to_unsigned(145, 8)),
			984 => std_logic_vector(to_unsigned(204, 8)),
			985 => std_logic_vector(to_unsigned(217, 8)),
			986 => std_logic_vector(to_unsigned(141, 8)),
			987 => std_logic_vector(to_unsigned(106, 8)),
			988 => std_logic_vector(to_unsigned(218, 8)),
			989 => std_logic_vector(to_unsigned(137, 8)),
			990 => std_logic_vector(to_unsigned(135, 8)),
			991 => std_logic_vector(to_unsigned(48, 8)),
			992 => std_logic_vector(to_unsigned(177, 8)),
			993 => std_logic_vector(to_unsigned(125, 8)),
			994 => std_logic_vector(to_unsigned(0, 8)),
			995 => std_logic_vector(to_unsigned(63, 8)),
			996 => std_logic_vector(to_unsigned(140, 8)),
			997 => std_logic_vector(to_unsigned(255, 8)),
			998 => std_logic_vector(to_unsigned(216, 8)),
			999 => std_logic_vector(to_unsigned(233, 8)),
			1000 => std_logic_vector(to_unsigned(157, 8)),
			1001 => std_logic_vector(to_unsigned(199, 8)),
			1002 => std_logic_vector(to_unsigned(232, 8)),
			1003 => std_logic_vector(to_unsigned(45, 8)),
			1004 => std_logic_vector(to_unsigned(86, 8)),
			1005 => std_logic_vector(to_unsigned(220, 8)),
			1006 => std_logic_vector(to_unsigned(79, 8)),
			1007 => std_logic_vector(to_unsigned(43, 8)),
			1008 => std_logic_vector(to_unsigned(226, 8)),
			1009 => std_logic_vector(to_unsigned(100, 8)),
			1010 => std_logic_vector(to_unsigned(158, 8)),
			1011 => std_logic_vector(to_unsigned(122, 8)),
			1012 => std_logic_vector(to_unsigned(28, 8)),
			1013 => std_logic_vector(to_unsigned(221, 8)),
			1014 => std_logic_vector(to_unsigned(2, 8)),
			1015 => std_logic_vector(to_unsigned(50, 8)),
			1016 => std_logic_vector(to_unsigned(159, 8)),
			1017 => std_logic_vector(to_unsigned(21, 8)),
			1018 => std_logic_vector(to_unsigned(245, 8)),
			1019 => std_logic_vector(to_unsigned(121, 8)),
			1020 => std_logic_vector(to_unsigned(237, 8)),
			1021 => std_logic_vector(to_unsigned(251, 8)),
			1022 => std_logic_vector(to_unsigned(106, 8)),
			1023 => std_logic_vector(to_unsigned(26, 8)),
			1024 => std_logic_vector(to_unsigned(243, 8)),
			1025 => std_logic_vector(to_unsigned(245, 8)),
			1026 => std_logic_vector(to_unsigned(253, 8)),
			1027 => std_logic_vector(to_unsigned(116, 8)),
			1028 => std_logic_vector(to_unsigned(205, 8)),
			1029 => std_logic_vector(to_unsigned(227, 8)),
			1030 => std_logic_vector(to_unsigned(94, 8)),
			1031 => std_logic_vector(to_unsigned(48, 8)),
			1032 => std_logic_vector(to_unsigned(90, 8)),
			1033 => std_logic_vector(to_unsigned(202, 8)),
			1034 => std_logic_vector(to_unsigned(78, 8)),
			1035 => std_logic_vector(to_unsigned(53, 8)),
			1036 => std_logic_vector(to_unsigned(74, 8)),
			1037 => std_logic_vector(to_unsigned(169, 8)),
			1038 => std_logic_vector(to_unsigned(186, 8)),
			1039 => std_logic_vector(to_unsigned(118, 8)),
			1040 => std_logic_vector(to_unsigned(249, 8)),
			1041 => std_logic_vector(to_unsigned(184, 8)),
			1042 => std_logic_vector(to_unsigned(59, 8)),
			1043 => std_logic_vector(to_unsigned(83, 8)),
			1044 => std_logic_vector(to_unsigned(21, 8)),
			1045 => std_logic_vector(to_unsigned(231, 8)),
			1046 => std_logic_vector(to_unsigned(132, 8)),
			1047 => std_logic_vector(to_unsigned(211, 8)),
			1048 => std_logic_vector(to_unsigned(203, 8)),
			1049 => std_logic_vector(to_unsigned(115, 8)),
			1050 => std_logic_vector(to_unsigned(108, 8)),
			1051 => std_logic_vector(to_unsigned(132, 8)),
			1052 => std_logic_vector(to_unsigned(183, 8)),
			1053 => std_logic_vector(to_unsigned(168, 8)),
			1054 => std_logic_vector(to_unsigned(75, 8)),
			1055 => std_logic_vector(to_unsigned(129, 8)),
			1056 => std_logic_vector(to_unsigned(121, 8)),
			1057 => std_logic_vector(to_unsigned(0, 8)),
			1058 => std_logic_vector(to_unsigned(119, 8)),
			1059 => std_logic_vector(to_unsigned(32, 8)),
			1060 => std_logic_vector(to_unsigned(145, 8)),
			1061 => std_logic_vector(to_unsigned(149, 8)),
			1062 => std_logic_vector(to_unsigned(107, 8)),
			1063 => std_logic_vector(to_unsigned(76, 8)),
			1064 => std_logic_vector(to_unsigned(84, 8)),
			1065 => std_logic_vector(to_unsigned(42, 8)),
			1066 => std_logic_vector(to_unsigned(178, 8)),
			1067 => std_logic_vector(to_unsigned(7, 8)),
			1068 => std_logic_vector(to_unsigned(196, 8)),
			1069 => std_logic_vector(to_unsigned(33, 8)),
			1070 => std_logic_vector(to_unsigned(159, 8)),
			1071 => std_logic_vector(to_unsigned(145, 8)),
			1072 => std_logic_vector(to_unsigned(169, 8)),
			1073 => std_logic_vector(to_unsigned(178, 8)),
			1074 => std_logic_vector(to_unsigned(136, 8)),
			1075 => std_logic_vector(to_unsigned(45, 8)),
			1076 => std_logic_vector(to_unsigned(14, 8)),
			1077 => std_logic_vector(to_unsigned(192, 8)),
			1078 => std_logic_vector(to_unsigned(43, 8)),
			1079 => std_logic_vector(to_unsigned(17, 8)),
			1080 => std_logic_vector(to_unsigned(71, 8)),
			1081 => std_logic_vector(to_unsigned(106, 8)),
			1082 => std_logic_vector(to_unsigned(3, 8)),
			1083 => std_logic_vector(to_unsigned(171, 8)),
			1084 => std_logic_vector(to_unsigned(244, 8)),
			1085 => std_logic_vector(to_unsigned(108, 8)),
			1086 => std_logic_vector(to_unsigned(166, 8)),
			1087 => std_logic_vector(to_unsigned(210, 8)),
			1088 => std_logic_vector(to_unsigned(148, 8)),
			1089 => std_logic_vector(to_unsigned(205, 8)),
			1090 => std_logic_vector(to_unsigned(164, 8)),
			1091 => std_logic_vector(to_unsigned(226, 8)),
			1092 => std_logic_vector(to_unsigned(204, 8)),
			1093 => std_logic_vector(to_unsigned(222, 8)),
			1094 => std_logic_vector(to_unsigned(145, 8)),
			1095 => std_logic_vector(to_unsigned(16, 8)),
			1096 => std_logic_vector(to_unsigned(211, 8)),
			1097 => std_logic_vector(to_unsigned(219, 8)),
			1098 => std_logic_vector(to_unsigned(70, 8)),
			1099 => std_logic_vector(to_unsigned(88, 8)),
			1100 => std_logic_vector(to_unsigned(173, 8)),
			1101 => std_logic_vector(to_unsigned(6, 8)),
			1102 => std_logic_vector(to_unsigned(39, 8)),
			1103 => std_logic_vector(to_unsigned(119, 8)),
			1104 => std_logic_vector(to_unsigned(164, 8)),
			1105 => std_logic_vector(to_unsigned(25, 8)),
			1106 => std_logic_vector(to_unsigned(4, 8)),
			1107 => std_logic_vector(to_unsigned(189, 8)),
			1108 => std_logic_vector(to_unsigned(32, 8)),
			1109 => std_logic_vector(to_unsigned(27, 8)),
			1110 => std_logic_vector(to_unsigned(173, 8)),
			1111 => std_logic_vector(to_unsigned(155, 8)),
			1112 => std_logic_vector(to_unsigned(110, 8)),
			1113 => std_logic_vector(to_unsigned(67, 8)),
			1114 => std_logic_vector(to_unsigned(85, 8)),
			1115 => std_logic_vector(to_unsigned(237, 8)),
			1116 => std_logic_vector(to_unsigned(164, 8)),
			1117 => std_logic_vector(to_unsigned(179, 8)),
			1118 => std_logic_vector(to_unsigned(117, 8)),
			1119 => std_logic_vector(to_unsigned(10, 8)),
			1120 => std_logic_vector(to_unsigned(217, 8)),
			1121 => std_logic_vector(to_unsigned(150, 8)),
			1122 => std_logic_vector(to_unsigned(144, 8)),
			1123 => std_logic_vector(to_unsigned(87, 8)),
			1124 => std_logic_vector(to_unsigned(208, 8)),
			1125 => std_logic_vector(to_unsigned(40, 8)),
			1126 => std_logic_vector(to_unsigned(167, 8)),
			1127 => std_logic_vector(to_unsigned(87, 8)),
			1128 => std_logic_vector(to_unsigned(242, 8)),
			1129 => std_logic_vector(to_unsigned(216, 8)),
			1130 => std_logic_vector(to_unsigned(111, 8)),
			1131 => std_logic_vector(to_unsigned(10, 8)),
			1132 => std_logic_vector(to_unsigned(43, 8)),
			1133 => std_logic_vector(to_unsigned(129, 8)),
			1134 => std_logic_vector(to_unsigned(178, 8)),
			1135 => std_logic_vector(to_unsigned(30, 8)),
			1136 => std_logic_vector(to_unsigned(130, 8)),
			1137 => std_logic_vector(to_unsigned(56, 8)),
			1138 => std_logic_vector(to_unsigned(143, 8)),
			1139 => std_logic_vector(to_unsigned(18, 8)),
			1140 => std_logic_vector(to_unsigned(143, 8)),
			1141 => std_logic_vector(to_unsigned(187, 8)),
			1142 => std_logic_vector(to_unsigned(247, 8)),
			1143 => std_logic_vector(to_unsigned(85, 8)),
			1144 => std_logic_vector(to_unsigned(147, 8)),
			1145 => std_logic_vector(to_unsigned(110, 8)),
			1146 => std_logic_vector(to_unsigned(244, 8)),
			1147 => std_logic_vector(to_unsigned(41, 8)),
			1148 => std_logic_vector(to_unsigned(46, 8)),
			1149 => std_logic_vector(to_unsigned(79, 8)),
			1150 => std_logic_vector(to_unsigned(182, 8)),
			1151 => std_logic_vector(to_unsigned(225, 8)),
			1152 => std_logic_vector(to_unsigned(255, 8)),
			1153 => std_logic_vector(to_unsigned(166, 8)),
			1154 => std_logic_vector(to_unsigned(190, 8)),
			1155 => std_logic_vector(to_unsigned(209, 8)),
			1156 => std_logic_vector(to_unsigned(163, 8)),
			1157 => std_logic_vector(to_unsigned(184, 8)),
			1158 => std_logic_vector(to_unsigned(11, 8)),
			1159 => std_logic_vector(to_unsigned(145, 8)),
			1160 => std_logic_vector(to_unsigned(112, 8)),
			1161 => std_logic_vector(to_unsigned(180, 8)),
			1162 => std_logic_vector(to_unsigned(201, 8)),
			1163 => std_logic_vector(to_unsigned(97, 8)),
			1164 => std_logic_vector(to_unsigned(84, 8)),
			1165 => std_logic_vector(to_unsigned(142, 8)),
			1166 => std_logic_vector(to_unsigned(244, 8)),
			1167 => std_logic_vector(to_unsigned(238, 8)),
			1168 => std_logic_vector(to_unsigned(156, 8)),
			1169 => std_logic_vector(to_unsigned(189, 8)),
			1170 => std_logic_vector(to_unsigned(65, 8)),
			1171 => std_logic_vector(to_unsigned(54, 8)),
			1172 => std_logic_vector(to_unsigned(178, 8)),
			1173 => std_logic_vector(to_unsigned(13, 8)),
			1174 => std_logic_vector(to_unsigned(108, 8)),
			1175 => std_logic_vector(to_unsigned(233, 8)),
			1176 => std_logic_vector(to_unsigned(105, 8)),
			1177 => std_logic_vector(to_unsigned(202, 8)),
			1178 => std_logic_vector(to_unsigned(163, 8)),
			1179 => std_logic_vector(to_unsigned(184, 8)),
			1180 => std_logic_vector(to_unsigned(217, 8)),
			1181 => std_logic_vector(to_unsigned(120, 8)),
			1182 => std_logic_vector(to_unsigned(69, 8)),
			1183 => std_logic_vector(to_unsigned(234, 8)),
			1184 => std_logic_vector(to_unsigned(66, 8)),
			1185 => std_logic_vector(to_unsigned(218, 8)),
			1186 => std_logic_vector(to_unsigned(63, 8)),
			1187 => std_logic_vector(to_unsigned(124, 8)),
			1188 => std_logic_vector(to_unsigned(242, 8)),
			1189 => std_logic_vector(to_unsigned(102, 8)),
			1190 => std_logic_vector(to_unsigned(47, 8)),
			1191 => std_logic_vector(to_unsigned(117, 8)),
			1192 => std_logic_vector(to_unsigned(161, 8)),
			1193 => std_logic_vector(to_unsigned(183, 8)),
			1194 => std_logic_vector(to_unsigned(181, 8)),
			1195 => std_logic_vector(to_unsigned(175, 8)),
			1196 => std_logic_vector(to_unsigned(182, 8)),
			1197 => std_logic_vector(to_unsigned(208, 8)),
			1198 => std_logic_vector(to_unsigned(158, 8)),
			1199 => std_logic_vector(to_unsigned(245, 8)),
			1200 => std_logic_vector(to_unsigned(96, 8)),
			1201 => std_logic_vector(to_unsigned(3, 8)),
			1202 => std_logic_vector(to_unsigned(161, 8)),
			1203 => std_logic_vector(to_unsigned(202, 8)),
			1204 => std_logic_vector(to_unsigned(8, 8)),
			1205 => std_logic_vector(to_unsigned(245, 8)),
			1206 => std_logic_vector(to_unsigned(71, 8)),
			1207 => std_logic_vector(to_unsigned(105, 8)),
			1208 => std_logic_vector(to_unsigned(217, 8)),
			1209 => std_logic_vector(to_unsigned(103, 8)),
			1210 => std_logic_vector(to_unsigned(198, 8)),
			1211 => std_logic_vector(to_unsigned(10, 8)),
			1212 => std_logic_vector(to_unsigned(10, 8)),
			1213 => std_logic_vector(to_unsigned(166, 8)),
			1214 => std_logic_vector(to_unsigned(100, 8)),
			1215 => std_logic_vector(to_unsigned(5, 8)),
			1216 => std_logic_vector(to_unsigned(109, 8)),
			1217 => std_logic_vector(to_unsigned(67, 8)),
			1218 => std_logic_vector(to_unsigned(86, 8)),
			1219 => std_logic_vector(to_unsigned(233, 8)),
			1220 => std_logic_vector(to_unsigned(145, 8)),
			1221 => std_logic_vector(to_unsigned(43, 8)),
			1222 => std_logic_vector(to_unsigned(74, 8)),
			1223 => std_logic_vector(to_unsigned(140, 8)),
			1224 => std_logic_vector(to_unsigned(115, 8)),
			1225 => std_logic_vector(to_unsigned(225, 8)),
			1226 => std_logic_vector(to_unsigned(222, 8)),
			1227 => std_logic_vector(to_unsigned(132, 8)),
			1228 => std_logic_vector(to_unsigned(199, 8)),
			1229 => std_logic_vector(to_unsigned(228, 8)),
			1230 => std_logic_vector(to_unsigned(182, 8)),
			1231 => std_logic_vector(to_unsigned(49, 8)),
			1232 => std_logic_vector(to_unsigned(196, 8)),
			1233 => std_logic_vector(to_unsigned(237, 8)),
			1234 => std_logic_vector(to_unsigned(202, 8)),
			1235 => std_logic_vector(to_unsigned(101, 8)),
			1236 => std_logic_vector(to_unsigned(235, 8)),
			1237 => std_logic_vector(to_unsigned(152, 8)),
			1238 => std_logic_vector(to_unsigned(71, 8)),
			1239 => std_logic_vector(to_unsigned(161, 8)),
			1240 => std_logic_vector(to_unsigned(244, 8)),
			1241 => std_logic_vector(to_unsigned(213, 8)),
			1242 => std_logic_vector(to_unsigned(168, 8)),
			1243 => std_logic_vector(to_unsigned(119, 8)),
			1244 => std_logic_vector(to_unsigned(160, 8)),
			1245 => std_logic_vector(to_unsigned(3, 8)),
			1246 => std_logic_vector(to_unsigned(128, 8)),
			1247 => std_logic_vector(to_unsigned(152, 8)),
			1248 => std_logic_vector(to_unsigned(231, 8)),
			1249 => std_logic_vector(to_unsigned(120, 8)),
			1250 => std_logic_vector(to_unsigned(58, 8)),
			1251 => std_logic_vector(to_unsigned(230, 8)),
			1252 => std_logic_vector(to_unsigned(52, 8)),
			1253 => std_logic_vector(to_unsigned(221, 8)),
			1254 => std_logic_vector(to_unsigned(167, 8)),
			1255 => std_logic_vector(to_unsigned(169, 8)),
			1256 => std_logic_vector(to_unsigned(23, 8)),
			1257 => std_logic_vector(to_unsigned(109, 8)),
			1258 => std_logic_vector(to_unsigned(35, 8)),
			1259 => std_logic_vector(to_unsigned(8, 8)),
			1260 => std_logic_vector(to_unsigned(212, 8)),
			1261 => std_logic_vector(to_unsigned(114, 8)),
			1262 => std_logic_vector(to_unsigned(224, 8)),
			1263 => std_logic_vector(to_unsigned(0, 8)),
			1264 => std_logic_vector(to_unsigned(228, 8)),
			1265 => std_logic_vector(to_unsigned(124, 8)),
			1266 => std_logic_vector(to_unsigned(166, 8)),
			1267 => std_logic_vector(to_unsigned(8, 8)),
			1268 => std_logic_vector(to_unsigned(72, 8)),
			1269 => std_logic_vector(to_unsigned(20, 8)),
			1270 => std_logic_vector(to_unsigned(211, 8)),
			1271 => std_logic_vector(to_unsigned(217, 8)),
			1272 => std_logic_vector(to_unsigned(173, 8)),
			1273 => std_logic_vector(to_unsigned(166, 8)),
			1274 => std_logic_vector(to_unsigned(230, 8)),
			1275 => std_logic_vector(to_unsigned(171, 8)),
			1276 => std_logic_vector(to_unsigned(50, 8)),
			1277 => std_logic_vector(to_unsigned(16, 8)),
			1278 => std_logic_vector(to_unsigned(22, 8)),
			1279 => std_logic_vector(to_unsigned(41, 8)),
			1280 => std_logic_vector(to_unsigned(131, 8)),
			1281 => std_logic_vector(to_unsigned(196, 8)),
			1282 => std_logic_vector(to_unsigned(161, 8)),
			1283 => std_logic_vector(to_unsigned(152, 8)),
			1284 => std_logic_vector(to_unsigned(132, 8)),
			1285 => std_logic_vector(to_unsigned(19, 8)),
			1286 => std_logic_vector(to_unsigned(82, 8)),
			1287 => std_logic_vector(to_unsigned(75, 8)),
			1288 => std_logic_vector(to_unsigned(141, 8)),
			1289 => std_logic_vector(to_unsigned(131, 8)),
			1290 => std_logic_vector(to_unsigned(230, 8)),
			1291 => std_logic_vector(to_unsigned(30, 8)),
			1292 => std_logic_vector(to_unsigned(232, 8)),
			1293 => std_logic_vector(to_unsigned(120, 8)),
			1294 => std_logic_vector(to_unsigned(203, 8)),
			1295 => std_logic_vector(to_unsigned(70, 8)),
			1296 => std_logic_vector(to_unsigned(122, 8)),
			1297 => std_logic_vector(to_unsigned(156, 8)),
			1298 => std_logic_vector(to_unsigned(143, 8)),
			1299 => std_logic_vector(to_unsigned(58, 8)),
			1300 => std_logic_vector(to_unsigned(225, 8)),
			1301 => std_logic_vector(to_unsigned(42, 8)),
			1302 => std_logic_vector(to_unsigned(194, 8)),
			1303 => std_logic_vector(to_unsigned(128, 8)),
			1304 => std_logic_vector(to_unsigned(164, 8)),
			1305 => std_logic_vector(to_unsigned(4, 8)),
			1306 => std_logic_vector(to_unsigned(131, 8)),
			1307 => std_logic_vector(to_unsigned(47, 8)),
			1308 => std_logic_vector(to_unsigned(125, 8)),
			1309 => std_logic_vector(to_unsigned(173, 8)),
			1310 => std_logic_vector(to_unsigned(43, 8)),
			1311 => std_logic_vector(to_unsigned(251, 8)),
			1312 => std_logic_vector(to_unsigned(246, 8)),
			1313 => std_logic_vector(to_unsigned(156, 8)),
			1314 => std_logic_vector(to_unsigned(162, 8)),
			1315 => std_logic_vector(to_unsigned(179, 8)),
			1316 => std_logic_vector(to_unsigned(217, 8)),
			1317 => std_logic_vector(to_unsigned(99, 8)),
			1318 => std_logic_vector(to_unsigned(146, 8)),
			1319 => std_logic_vector(to_unsigned(114, 8)),
			1320 => std_logic_vector(to_unsigned(79, 8)),
			1321 => std_logic_vector(to_unsigned(39, 8)),
			1322 => std_logic_vector(to_unsigned(151, 8)),
			1323 => std_logic_vector(to_unsigned(140, 8)),
			1324 => std_logic_vector(to_unsigned(232, 8)),
			1325 => std_logic_vector(to_unsigned(201, 8)),
			1326 => std_logic_vector(to_unsigned(114, 8)),
			1327 => std_logic_vector(to_unsigned(106, 8)),
			1328 => std_logic_vector(to_unsigned(200, 8)),
			1329 => std_logic_vector(to_unsigned(17, 8)),
			1330 => std_logic_vector(to_unsigned(210, 8)),
			1331 => std_logic_vector(to_unsigned(237, 8)),
			1332 => std_logic_vector(to_unsigned(48, 8)),
			1333 => std_logic_vector(to_unsigned(81, 8)),
			1334 => std_logic_vector(to_unsigned(216, 8)),
			1335 => std_logic_vector(to_unsigned(207, 8)),
			1336 => std_logic_vector(to_unsigned(249, 8)),
			1337 => std_logic_vector(to_unsigned(220, 8)),
			1338 => std_logic_vector(to_unsigned(205, 8)),
			1339 => std_logic_vector(to_unsigned(212, 8)),
			1340 => std_logic_vector(to_unsigned(211, 8)),
			1341 => std_logic_vector(to_unsigned(75, 8)),
			1342 => std_logic_vector(to_unsigned(111, 8)),
			1343 => std_logic_vector(to_unsigned(184, 8)),
			1344 => std_logic_vector(to_unsigned(60, 8)),
			1345 => std_logic_vector(to_unsigned(204, 8)),
			1346 => std_logic_vector(to_unsigned(52, 8)),
			1347 => std_logic_vector(to_unsigned(201, 8)),
			1348 => std_logic_vector(to_unsigned(186, 8)),
			1349 => std_logic_vector(to_unsigned(108, 8)),
			1350 => std_logic_vector(to_unsigned(91, 8)),
			1351 => std_logic_vector(to_unsigned(205, 8)),
			1352 => std_logic_vector(to_unsigned(65, 8)),
			1353 => std_logic_vector(to_unsigned(129, 8)),
			1354 => std_logic_vector(to_unsigned(216, 8)),
			1355 => std_logic_vector(to_unsigned(244, 8)),
			1356 => std_logic_vector(to_unsigned(238, 8)),
			1357 => std_logic_vector(to_unsigned(86, 8)),
			1358 => std_logic_vector(to_unsigned(179, 8)),
			1359 => std_logic_vector(to_unsigned(76, 8)),
			1360 => std_logic_vector(to_unsigned(248, 8)),
			1361 => std_logic_vector(to_unsigned(141, 8)),
			1362 => std_logic_vector(to_unsigned(197, 8)),
			1363 => std_logic_vector(to_unsigned(207, 8)),
			1364 => std_logic_vector(to_unsigned(68, 8)),
			1365 => std_logic_vector(to_unsigned(114, 8)),
			1366 => std_logic_vector(to_unsigned(68, 8)),
			1367 => std_logic_vector(to_unsigned(82, 8)),
			1368 => std_logic_vector(to_unsigned(76, 8)),
			1369 => std_logic_vector(to_unsigned(82, 8)),
			1370 => std_logic_vector(to_unsigned(14, 8)),
			1371 => std_logic_vector(to_unsigned(119, 8)),
			1372 => std_logic_vector(to_unsigned(165, 8)),
			1373 => std_logic_vector(to_unsigned(211, 8)),
			1374 => std_logic_vector(to_unsigned(127, 8)),
			1375 => std_logic_vector(to_unsigned(68, 8)),
			1376 => std_logic_vector(to_unsigned(231, 8)),
			1377 => std_logic_vector(to_unsigned(174, 8)),
			1378 => std_logic_vector(to_unsigned(164, 8)),
			1379 => std_logic_vector(to_unsigned(65, 8)),
			1380 => std_logic_vector(to_unsigned(63, 8)),
			1381 => std_logic_vector(to_unsigned(0, 8)),
			1382 => std_logic_vector(to_unsigned(35, 8)),
			1383 => std_logic_vector(to_unsigned(92, 8)),
			1384 => std_logic_vector(to_unsigned(75, 8)),
			1385 => std_logic_vector(to_unsigned(96, 8)),
			1386 => std_logic_vector(to_unsigned(1, 8)),
			1387 => std_logic_vector(to_unsigned(203, 8)),
			1388 => std_logic_vector(to_unsigned(254, 8)),
			1389 => std_logic_vector(to_unsigned(219, 8)),
			1390 => std_logic_vector(to_unsigned(222, 8)),
			1391 => std_logic_vector(to_unsigned(248, 8)),
			1392 => std_logic_vector(to_unsigned(168, 8)),
			1393 => std_logic_vector(to_unsigned(186, 8)),
			1394 => std_logic_vector(to_unsigned(241, 8)),
			1395 => std_logic_vector(to_unsigned(185, 8)),
			1396 => std_logic_vector(to_unsigned(117, 8)),
			1397 => std_logic_vector(to_unsigned(128, 8)),
			1398 => std_logic_vector(to_unsigned(243, 8)),
			1399 => std_logic_vector(to_unsigned(44, 8)),
			1400 => std_logic_vector(to_unsigned(222, 8)),
			1401 => std_logic_vector(to_unsigned(168, 8)),
			1402 => std_logic_vector(to_unsigned(222, 8)),
			1403 => std_logic_vector(to_unsigned(161, 8)),
			1404 => std_logic_vector(to_unsigned(51, 8)),
			1405 => std_logic_vector(to_unsigned(14, 8)),
			1406 => std_logic_vector(to_unsigned(107, 8)),
			1407 => std_logic_vector(to_unsigned(68, 8)),
			1408 => std_logic_vector(to_unsigned(74, 8)),
			1409 => std_logic_vector(to_unsigned(106, 8)),
			1410 => std_logic_vector(to_unsigned(0, 8)),
			1411 => std_logic_vector(to_unsigned(45, 8)),
			1412 => std_logic_vector(to_unsigned(223, 8)),
			1413 => std_logic_vector(to_unsigned(0, 8)),
			1414 => std_logic_vector(to_unsigned(201, 8)),
			1415 => std_logic_vector(to_unsigned(28, 8)),
			1416 => std_logic_vector(to_unsigned(221, 8)),
			1417 => std_logic_vector(to_unsigned(92, 8)),
			1418 => std_logic_vector(to_unsigned(151, 8)),
			1419 => std_logic_vector(to_unsigned(112, 8)),
			1420 => std_logic_vector(to_unsigned(130, 8)),
			1421 => std_logic_vector(to_unsigned(234, 8)),
			1422 => std_logic_vector(to_unsigned(89, 8)),
			1423 => std_logic_vector(to_unsigned(47, 8)),
			1424 => std_logic_vector(to_unsigned(103, 8)),
			1425 => std_logic_vector(to_unsigned(46, 8)),
			1426 => std_logic_vector(to_unsigned(73, 8)),
			1427 => std_logic_vector(to_unsigned(123, 8)),
			1428 => std_logic_vector(to_unsigned(31, 8)),
			1429 => std_logic_vector(to_unsigned(9, 8)),
			1430 => std_logic_vector(to_unsigned(31, 8)),
			1431 => std_logic_vector(to_unsigned(45, 8)),
			1432 => std_logic_vector(to_unsigned(66, 8)),
			1433 => std_logic_vector(to_unsigned(55, 8)),
			1434 => std_logic_vector(to_unsigned(103, 8)),
			1435 => std_logic_vector(to_unsigned(166, 8)),
			1436 => std_logic_vector(to_unsigned(110, 8)),
			1437 => std_logic_vector(to_unsigned(233, 8)),
			1438 => std_logic_vector(to_unsigned(108, 8)),
			1439 => std_logic_vector(to_unsigned(111, 8)),
			1440 => std_logic_vector(to_unsigned(41, 8)),
			1441 => std_logic_vector(to_unsigned(148, 8)),
			1442 => std_logic_vector(to_unsigned(194, 8)),
			1443 => std_logic_vector(to_unsigned(99, 8)),
			1444 => std_logic_vector(to_unsigned(116, 8)),
			1445 => std_logic_vector(to_unsigned(166, 8)),
			1446 => std_logic_vector(to_unsigned(185, 8)),
			1447 => std_logic_vector(to_unsigned(144, 8)),
			1448 => std_logic_vector(to_unsigned(192, 8)),
			1449 => std_logic_vector(to_unsigned(214, 8)),
			1450 => std_logic_vector(to_unsigned(78, 8)),
			1451 => std_logic_vector(to_unsigned(90, 8)),
			1452 => std_logic_vector(to_unsigned(20, 8)),
			1453 => std_logic_vector(to_unsigned(132, 8)),
			1454 => std_logic_vector(to_unsigned(79, 8)),
			1455 => std_logic_vector(to_unsigned(29, 8)),
			1456 => std_logic_vector(to_unsigned(12, 8)),
			1457 => std_logic_vector(to_unsigned(86, 8)),
			1458 => std_logic_vector(to_unsigned(58, 8)),
			1459 => std_logic_vector(to_unsigned(168, 8)),
			1460 => std_logic_vector(to_unsigned(127, 8)),
			1461 => std_logic_vector(to_unsigned(133, 8)),
			1462 => std_logic_vector(to_unsigned(1, 8)),
			1463 => std_logic_vector(to_unsigned(49, 8)),
			1464 => std_logic_vector(to_unsigned(26, 8)),
			1465 => std_logic_vector(to_unsigned(126, 8)),
			1466 => std_logic_vector(to_unsigned(151, 8)),
			1467 => std_logic_vector(to_unsigned(5, 8)),
			1468 => std_logic_vector(to_unsigned(225, 8)),
			1469 => std_logic_vector(to_unsigned(47, 8)),
			1470 => std_logic_vector(to_unsigned(131, 8)),
			1471 => std_logic_vector(to_unsigned(73, 8)),
			1472 => std_logic_vector(to_unsigned(78, 8)),
			1473 => std_logic_vector(to_unsigned(163, 8)),
			1474 => std_logic_vector(to_unsigned(85, 8)),
			1475 => std_logic_vector(to_unsigned(191, 8)),
			1476 => std_logic_vector(to_unsigned(32, 8)),
			1477 => std_logic_vector(to_unsigned(70, 8)),
			1478 => std_logic_vector(to_unsigned(228, 8)),
			1479 => std_logic_vector(to_unsigned(133, 8)),
			1480 => std_logic_vector(to_unsigned(208, 8)),
			1481 => std_logic_vector(to_unsigned(105, 8)),
			1482 => std_logic_vector(to_unsigned(39, 8)),
			1483 => std_logic_vector(to_unsigned(39, 8)),
			1484 => std_logic_vector(to_unsigned(64, 8)),
			1485 => std_logic_vector(to_unsigned(238, 8)),
			1486 => std_logic_vector(to_unsigned(146, 8)),
			1487 => std_logic_vector(to_unsigned(5, 8)),
			1488 => std_logic_vector(to_unsigned(227, 8)),
			1489 => std_logic_vector(to_unsigned(177, 8)),
			1490 => std_logic_vector(to_unsigned(210, 8)),
			1491 => std_logic_vector(to_unsigned(237, 8)),
			1492 => std_logic_vector(to_unsigned(182, 8)),
			1493 => std_logic_vector(to_unsigned(231, 8)),
			1494 => std_logic_vector(to_unsigned(241, 8)),
			1495 => std_logic_vector(to_unsigned(188, 8)),
			1496 => std_logic_vector(to_unsigned(46, 8)),
			1497 => std_logic_vector(to_unsigned(57, 8)),
			1498 => std_logic_vector(to_unsigned(239, 8)),
			1499 => std_logic_vector(to_unsigned(101, 8)),
			1500 => std_logic_vector(to_unsigned(221, 8)),
			1501 => std_logic_vector(to_unsigned(41, 8)),
			1502 => std_logic_vector(to_unsigned(112, 8)),
			1503 => std_logic_vector(to_unsigned(157, 8)),
			1504 => std_logic_vector(to_unsigned(207, 8)),
			1505 => std_logic_vector(to_unsigned(81, 8)),
			1506 => std_logic_vector(to_unsigned(201, 8)),
			1507 => std_logic_vector(to_unsigned(233, 8)),
			1508 => std_logic_vector(to_unsigned(116, 8)),
			1509 => std_logic_vector(to_unsigned(82, 8)),
			1510 => std_logic_vector(to_unsigned(49, 8)),
			1511 => std_logic_vector(to_unsigned(2, 8)),
			1512 => std_logic_vector(to_unsigned(194, 8)),
			1513 => std_logic_vector(to_unsigned(151, 8)),
			1514 => std_logic_vector(to_unsigned(8, 8)),
			1515 => std_logic_vector(to_unsigned(162, 8)),
			1516 => std_logic_vector(to_unsigned(198, 8)),
			1517 => std_logic_vector(to_unsigned(246, 8)),
			1518 => std_logic_vector(to_unsigned(111, 8)),
			1519 => std_logic_vector(to_unsigned(220, 8)),
			1520 => std_logic_vector(to_unsigned(100, 8)),
			1521 => std_logic_vector(to_unsigned(90, 8)),
			1522 => std_logic_vector(to_unsigned(216, 8)),
			1523 => std_logic_vector(to_unsigned(205, 8)),
			1524 => std_logic_vector(to_unsigned(174, 8)),
			1525 => std_logic_vector(to_unsigned(85, 8)),
			1526 => std_logic_vector(to_unsigned(107, 8)),
			1527 => std_logic_vector(to_unsigned(19, 8)),
			1528 => std_logic_vector(to_unsigned(24, 8)),
			1529 => std_logic_vector(to_unsigned(73, 8)),
			1530 => std_logic_vector(to_unsigned(23, 8)),
			1531 => std_logic_vector(to_unsigned(189, 8)),
			1532 => std_logic_vector(to_unsigned(205, 8)),
			1533 => std_logic_vector(to_unsigned(120, 8)),
			1534 => std_logic_vector(to_unsigned(134, 8)),
			1535 => std_logic_vector(to_unsigned(219, 8)),
			1536 => std_logic_vector(to_unsigned(16, 8)),
			1537 => std_logic_vector(to_unsigned(142, 8)),
			1538 => std_logic_vector(to_unsigned(239, 8)),
			1539 => std_logic_vector(to_unsigned(122, 8)),
			1540 => std_logic_vector(to_unsigned(122, 8)),
			1541 => std_logic_vector(to_unsigned(47, 8)),
			1542 => std_logic_vector(to_unsigned(73, 8)),
			1543 => std_logic_vector(to_unsigned(83, 8)),
			1544 => std_logic_vector(to_unsigned(155, 8)),
			1545 => std_logic_vector(to_unsigned(235, 8)),
			1546 => std_logic_vector(to_unsigned(155, 8)),
			1547 => std_logic_vector(to_unsigned(153, 8)),
			1548 => std_logic_vector(to_unsigned(50, 8)),
			1549 => std_logic_vector(to_unsigned(216, 8)),
			1550 => std_logic_vector(to_unsigned(233, 8)),
			1551 => std_logic_vector(to_unsigned(66, 8)),
			1552 => std_logic_vector(to_unsigned(88, 8)),
			1553 => std_logic_vector(to_unsigned(79, 8)),
			1554 => std_logic_vector(to_unsigned(196, 8)),
			1555 => std_logic_vector(to_unsigned(64, 8)),
			1556 => std_logic_vector(to_unsigned(156, 8)),
			1557 => std_logic_vector(to_unsigned(25, 8)),
			1558 => std_logic_vector(to_unsigned(184, 8)),
			1559 => std_logic_vector(to_unsigned(108, 8)),
			1560 => std_logic_vector(to_unsigned(155, 8)),
			1561 => std_logic_vector(to_unsigned(74, 8)),
			1562 => std_logic_vector(to_unsigned(205, 8)),
			1563 => std_logic_vector(to_unsigned(10, 8)),
			1564 => std_logic_vector(to_unsigned(228, 8)),
			1565 => std_logic_vector(to_unsigned(87, 8)),
			1566 => std_logic_vector(to_unsigned(7, 8)),
			1567 => std_logic_vector(to_unsigned(145, 8)),
			1568 => std_logic_vector(to_unsigned(18, 8)),
			1569 => std_logic_vector(to_unsigned(59, 8)),
			1570 => std_logic_vector(to_unsigned(71, 8)),
			1571 => std_logic_vector(to_unsigned(91, 8)),
			1572 => std_logic_vector(to_unsigned(75, 8)),
			1573 => std_logic_vector(to_unsigned(179, 8)),
			1574 => std_logic_vector(to_unsigned(232, 8)),
			1575 => std_logic_vector(to_unsigned(23, 8)),
			1576 => std_logic_vector(to_unsigned(20, 8)),
			1577 => std_logic_vector(to_unsigned(79, 8)),
			1578 => std_logic_vector(to_unsigned(183, 8)),
			1579 => std_logic_vector(to_unsigned(67, 8)),
			1580 => std_logic_vector(to_unsigned(185, 8)),
			1581 => std_logic_vector(to_unsigned(13, 8)),
			1582 => std_logic_vector(to_unsigned(38, 8)),
			1583 => std_logic_vector(to_unsigned(52, 8)),
			1584 => std_logic_vector(to_unsigned(134, 8)),
			1585 => std_logic_vector(to_unsigned(210, 8)),
			1586 => std_logic_vector(to_unsigned(165, 8)),
			1587 => std_logic_vector(to_unsigned(235, 8)),
			1588 => std_logic_vector(to_unsigned(162, 8)),
			1589 => std_logic_vector(to_unsigned(201, 8)),
			1590 => std_logic_vector(to_unsigned(18, 8)),
			1591 => std_logic_vector(to_unsigned(198, 8)),
			1592 => std_logic_vector(to_unsigned(7, 8)),
			1593 => std_logic_vector(to_unsigned(42, 8)),
			1594 => std_logic_vector(to_unsigned(191, 8)),
			1595 => std_logic_vector(to_unsigned(89, 8)),
			1596 => std_logic_vector(to_unsigned(162, 8)),
			1597 => std_logic_vector(to_unsigned(216, 8)),
			1598 => std_logic_vector(to_unsigned(34, 8)),
			1599 => std_logic_vector(to_unsigned(164, 8)),
			1600 => std_logic_vector(to_unsigned(180, 8)),
			1601 => std_logic_vector(to_unsigned(188, 8)),
			1602 => std_logic_vector(to_unsigned(250, 8)),
			1603 => std_logic_vector(to_unsigned(27, 8)),
			1604 => std_logic_vector(to_unsigned(190, 8)),
			1605 => std_logic_vector(to_unsigned(114, 8)),
			1606 => std_logic_vector(to_unsigned(183, 8)),
			1607 => std_logic_vector(to_unsigned(248, 8)),
			1608 => std_logic_vector(to_unsigned(203, 8)),
			1609 => std_logic_vector(to_unsigned(24, 8)),
			1610 => std_logic_vector(to_unsigned(179, 8)),
			1611 => std_logic_vector(to_unsigned(75, 8)),
			1612 => std_logic_vector(to_unsigned(11, 8)),
			1613 => std_logic_vector(to_unsigned(123, 8)),
			1614 => std_logic_vector(to_unsigned(97, 8)),
			1615 => std_logic_vector(to_unsigned(27, 8)),
			1616 => std_logic_vector(to_unsigned(177, 8)),
			1617 => std_logic_vector(to_unsigned(112, 8)),
			1618 => std_logic_vector(to_unsigned(17, 8)),
			1619 => std_logic_vector(to_unsigned(126, 8)),
			1620 => std_logic_vector(to_unsigned(37, 8)),
			1621 => std_logic_vector(to_unsigned(227, 8)),
			1622 => std_logic_vector(to_unsigned(11, 8)),
			1623 => std_logic_vector(to_unsigned(131, 8)),
			1624 => std_logic_vector(to_unsigned(119, 8)),
			1625 => std_logic_vector(to_unsigned(31, 8)),
			1626 => std_logic_vector(to_unsigned(50, 8)),
			1627 => std_logic_vector(to_unsigned(37, 8)),
			1628 => std_logic_vector(to_unsigned(117, 8)),
			1629 => std_logic_vector(to_unsigned(203, 8)),
			1630 => std_logic_vector(to_unsigned(235, 8)),
			1631 => std_logic_vector(to_unsigned(27, 8)),
			1632 => std_logic_vector(to_unsigned(4, 8)),
			1633 => std_logic_vector(to_unsigned(124, 8)),
			1634 => std_logic_vector(to_unsigned(190, 8)),
			1635 => std_logic_vector(to_unsigned(24, 8)),
			1636 => std_logic_vector(to_unsigned(38, 8)),
			1637 => std_logic_vector(to_unsigned(105, 8)),
			1638 => std_logic_vector(to_unsigned(182, 8)),
			1639 => std_logic_vector(to_unsigned(130, 8)),
			1640 => std_logic_vector(to_unsigned(209, 8)),
			1641 => std_logic_vector(to_unsigned(191, 8)),
			1642 => std_logic_vector(to_unsigned(13, 8)),
			1643 => std_logic_vector(to_unsigned(41, 8)),
			1644 => std_logic_vector(to_unsigned(235, 8)),
			1645 => std_logic_vector(to_unsigned(114, 8)),
			1646 => std_logic_vector(to_unsigned(28, 8)),
			1647 => std_logic_vector(to_unsigned(192, 8)),
			1648 => std_logic_vector(to_unsigned(9, 8)),
			1649 => std_logic_vector(to_unsigned(144, 8)),
			1650 => std_logic_vector(to_unsigned(61, 8)),
			1651 => std_logic_vector(to_unsigned(93, 8)),
			1652 => std_logic_vector(to_unsigned(85, 8)),
			1653 => std_logic_vector(to_unsigned(9, 8)),
			1654 => std_logic_vector(to_unsigned(246, 8)),
			1655 => std_logic_vector(to_unsigned(144, 8)),
			1656 => std_logic_vector(to_unsigned(177, 8)),
			1657 => std_logic_vector(to_unsigned(65, 8)),
			1658 => std_logic_vector(to_unsigned(68, 8)),
			1659 => std_logic_vector(to_unsigned(48, 8)),
			1660 => std_logic_vector(to_unsigned(180, 8)),
			1661 => std_logic_vector(to_unsigned(129, 8)),
			1662 => std_logic_vector(to_unsigned(129, 8)),
			1663 => std_logic_vector(to_unsigned(244, 8)),
			1664 => std_logic_vector(to_unsigned(220, 8)),
			1665 => std_logic_vector(to_unsigned(63, 8)),
			1666 => std_logic_vector(to_unsigned(3, 8)),
			1667 => std_logic_vector(to_unsigned(244, 8)),
			1668 => std_logic_vector(to_unsigned(44, 8)),
			1669 => std_logic_vector(to_unsigned(19, 8)),
			1670 => std_logic_vector(to_unsigned(79, 8)),
			1671 => std_logic_vector(to_unsigned(81, 8)),
			1672 => std_logic_vector(to_unsigned(148, 8)),
			1673 => std_logic_vector(to_unsigned(154, 8)),
			1674 => std_logic_vector(to_unsigned(158, 8)),
			1675 => std_logic_vector(to_unsigned(52, 8)),
			1676 => std_logic_vector(to_unsigned(136, 8)),
			1677 => std_logic_vector(to_unsigned(121, 8)),
			1678 => std_logic_vector(to_unsigned(230, 8)),
			1679 => std_logic_vector(to_unsigned(31, 8)),
			1680 => std_logic_vector(to_unsigned(171, 8)),
			1681 => std_logic_vector(to_unsigned(2, 8)),
			1682 => std_logic_vector(to_unsigned(49, 8)),
			1683 => std_logic_vector(to_unsigned(23, 8)),
			1684 => std_logic_vector(to_unsigned(125, 8)),
			1685 => std_logic_vector(to_unsigned(255, 8)),
			1686 => std_logic_vector(to_unsigned(175, 8)),
			1687 => std_logic_vector(to_unsigned(246, 8)),
			1688 => std_logic_vector(to_unsigned(57, 8)),
			1689 => std_logic_vector(to_unsigned(23, 8)),
			1690 => std_logic_vector(to_unsigned(221, 8)),
			1691 => std_logic_vector(to_unsigned(138, 8)),
			1692 => std_logic_vector(to_unsigned(181, 8)),
			1693 => std_logic_vector(to_unsigned(189, 8)),
			1694 => std_logic_vector(to_unsigned(28, 8)),
			1695 => std_logic_vector(to_unsigned(16, 8)),
			1696 => std_logic_vector(to_unsigned(193, 8)),
			1697 => std_logic_vector(to_unsigned(30, 8)),
			1698 => std_logic_vector(to_unsigned(179, 8)),
			1699 => std_logic_vector(to_unsigned(222, 8)),
			1700 => std_logic_vector(to_unsigned(78, 8)),
			1701 => std_logic_vector(to_unsigned(243, 8)),
			1702 => std_logic_vector(to_unsigned(16, 8)),
			1703 => std_logic_vector(to_unsigned(142, 8)),
			1704 => std_logic_vector(to_unsigned(232, 8)),
			1705 => std_logic_vector(to_unsigned(248, 8)),
			1706 => std_logic_vector(to_unsigned(88, 8)),
			1707 => std_logic_vector(to_unsigned(175, 8)),
			1708 => std_logic_vector(to_unsigned(101, 8)),
			1709 => std_logic_vector(to_unsigned(130, 8)),
			1710 => std_logic_vector(to_unsigned(91, 8)),
			1711 => std_logic_vector(to_unsigned(7, 8)),
			1712 => std_logic_vector(to_unsigned(197, 8)),
			1713 => std_logic_vector(to_unsigned(138, 8)),
			1714 => std_logic_vector(to_unsigned(129, 8)),
			1715 => std_logic_vector(to_unsigned(228, 8)),
			1716 => std_logic_vector(to_unsigned(187, 8)),
			1717 => std_logic_vector(to_unsigned(106, 8)),
			1718 => std_logic_vector(to_unsigned(186, 8)),
			1719 => std_logic_vector(to_unsigned(80, 8)),
			1720 => std_logic_vector(to_unsigned(93, 8)),
			1721 => std_logic_vector(to_unsigned(38, 8)),
			1722 => std_logic_vector(to_unsigned(13, 8)),
			1723 => std_logic_vector(to_unsigned(29, 8)),
			1724 => std_logic_vector(to_unsigned(90, 8)),
			1725 => std_logic_vector(to_unsigned(7, 8)),
			1726 => std_logic_vector(to_unsigned(70, 8)),
			1727 => std_logic_vector(to_unsigned(143, 8)),
			1728 => std_logic_vector(to_unsigned(226, 8)),
			1729 => std_logic_vector(to_unsigned(83, 8)),
			1730 => std_logic_vector(to_unsigned(246, 8)),
			1731 => std_logic_vector(to_unsigned(71, 8)),
			1732 => std_logic_vector(to_unsigned(241, 8)),
			1733 => std_logic_vector(to_unsigned(210, 8)),
			1734 => std_logic_vector(to_unsigned(116, 8)),
			1735 => std_logic_vector(to_unsigned(99, 8)),
			1736 => std_logic_vector(to_unsigned(137, 8)),
			1737 => std_logic_vector(to_unsigned(29, 8)),
			1738 => std_logic_vector(to_unsigned(54, 8)),
			1739 => std_logic_vector(to_unsigned(105, 8)),
			1740 => std_logic_vector(to_unsigned(168, 8)),
			1741 => std_logic_vector(to_unsigned(67, 8)),
			1742 => std_logic_vector(to_unsigned(240, 8)),
			1743 => std_logic_vector(to_unsigned(55, 8)),
			1744 => std_logic_vector(to_unsigned(235, 8)),
			1745 => std_logic_vector(to_unsigned(204, 8)),
			1746 => std_logic_vector(to_unsigned(109, 8)),
			1747 => std_logic_vector(to_unsigned(51, 8)),
			1748 => std_logic_vector(to_unsigned(228, 8)),
			1749 => std_logic_vector(to_unsigned(110, 8)),
			1750 => std_logic_vector(to_unsigned(156, 8)),
			1751 => std_logic_vector(to_unsigned(69, 8)),
			1752 => std_logic_vector(to_unsigned(177, 8)),
			1753 => std_logic_vector(to_unsigned(13, 8)),
			1754 => std_logic_vector(to_unsigned(197, 8)),
			1755 => std_logic_vector(to_unsigned(190, 8)),
			1756 => std_logic_vector(to_unsigned(150, 8)),
			1757 => std_logic_vector(to_unsigned(28, 8)),
			1758 => std_logic_vector(to_unsigned(114, 8)),
			1759 => std_logic_vector(to_unsigned(211, 8)),
			1760 => std_logic_vector(to_unsigned(193, 8)),
			1761 => std_logic_vector(to_unsigned(228, 8)),
			1762 => std_logic_vector(to_unsigned(131, 8)),
			1763 => std_logic_vector(to_unsigned(210, 8)),
			1764 => std_logic_vector(to_unsigned(248, 8)),
			1765 => std_logic_vector(to_unsigned(66, 8)),
			1766 => std_logic_vector(to_unsigned(140, 8)),
			1767 => std_logic_vector(to_unsigned(119, 8)),
			1768 => std_logic_vector(to_unsigned(115, 8)),
			1769 => std_logic_vector(to_unsigned(179, 8)),
			1770 => std_logic_vector(to_unsigned(32, 8)),
			1771 => std_logic_vector(to_unsigned(71, 8)),
			1772 => std_logic_vector(to_unsigned(1, 8)),
			1773 => std_logic_vector(to_unsigned(55, 8)),
			1774 => std_logic_vector(to_unsigned(108, 8)),
			1775 => std_logic_vector(to_unsigned(87, 8)),
			1776 => std_logic_vector(to_unsigned(187, 8)),
			1777 => std_logic_vector(to_unsigned(29, 8)),
			1778 => std_logic_vector(to_unsigned(252, 8)),
			1779 => std_logic_vector(to_unsigned(140, 8)),
			1780 => std_logic_vector(to_unsigned(212, 8)),
			1781 => std_logic_vector(to_unsigned(247, 8)),
			1782 => std_logic_vector(to_unsigned(129, 8)),
			1783 => std_logic_vector(to_unsigned(230, 8)),
			1784 => std_logic_vector(to_unsigned(5, 8)),
			1785 => std_logic_vector(to_unsigned(201, 8)),
			1786 => std_logic_vector(to_unsigned(254, 8)),
			1787 => std_logic_vector(to_unsigned(59, 8)),
			1788 => std_logic_vector(to_unsigned(208, 8)),
			1789 => std_logic_vector(to_unsigned(226, 8)),
			1790 => std_logic_vector(to_unsigned(123, 8)),
			1791 => std_logic_vector(to_unsigned(127, 8)),
			1792 => std_logic_vector(to_unsigned(255, 8)),
			1793 => std_logic_vector(to_unsigned(13, 8)),
			1794 => std_logic_vector(to_unsigned(246, 8)),
			1795 => std_logic_vector(to_unsigned(126, 8)),
			1796 => std_logic_vector(to_unsigned(233, 8)),
			1797 => std_logic_vector(to_unsigned(189, 8)),
			1798 => std_logic_vector(to_unsigned(136, 8)),
			1799 => std_logic_vector(to_unsigned(58, 8)),
			1800 => std_logic_vector(to_unsigned(160, 8)),
			1801 => std_logic_vector(to_unsigned(145, 8)),
			1802 => std_logic_vector(to_unsigned(64, 8)),
			1803 => std_logic_vector(to_unsigned(72, 8)),
			1804 => std_logic_vector(to_unsigned(229, 8)),
			1805 => std_logic_vector(to_unsigned(123, 8)),
			1806 => std_logic_vector(to_unsigned(177, 8)),
			1807 => std_logic_vector(to_unsigned(201, 8)),
			1808 => std_logic_vector(to_unsigned(8, 8)),
			1809 => std_logic_vector(to_unsigned(179, 8)),
			1810 => std_logic_vector(to_unsigned(237, 8)),
			1811 => std_logic_vector(to_unsigned(248, 8)),
			1812 => std_logic_vector(to_unsigned(151, 8)),
			1813 => std_logic_vector(to_unsigned(215, 8)),
			1814 => std_logic_vector(to_unsigned(74, 8)),
			1815 => std_logic_vector(to_unsigned(48, 8)),
			1816 => std_logic_vector(to_unsigned(90, 8)),
			1817 => std_logic_vector(to_unsigned(64, 8)),
			1818 => std_logic_vector(to_unsigned(185, 8)),
			1819 => std_logic_vector(to_unsigned(67, 8)),
			1820 => std_logic_vector(to_unsigned(21, 8)),
			1821 => std_logic_vector(to_unsigned(166, 8)),
			1822 => std_logic_vector(to_unsigned(103, 8)),
			1823 => std_logic_vector(to_unsigned(22, 8)),
			1824 => std_logic_vector(to_unsigned(190, 8)),
			1825 => std_logic_vector(to_unsigned(172, 8)),
			1826 => std_logic_vector(to_unsigned(83, 8)),
			1827 => std_logic_vector(to_unsigned(207, 8)),
			1828 => std_logic_vector(to_unsigned(77, 8)),
			1829 => std_logic_vector(to_unsigned(3, 8)),
			1830 => std_logic_vector(to_unsigned(64, 8)),
			1831 => std_logic_vector(to_unsigned(182, 8)),
			1832 => std_logic_vector(to_unsigned(152, 8)),
			1833 => std_logic_vector(to_unsigned(11, 8)),
			1834 => std_logic_vector(to_unsigned(76, 8)),
			1835 => std_logic_vector(to_unsigned(47, 8)),
			1836 => std_logic_vector(to_unsigned(79, 8)),
			1837 => std_logic_vector(to_unsigned(97, 8)),
			1838 => std_logic_vector(to_unsigned(200, 8)),
			1839 => std_logic_vector(to_unsigned(35, 8)),
			1840 => std_logic_vector(to_unsigned(203, 8)),
			1841 => std_logic_vector(to_unsigned(187, 8)),
			1842 => std_logic_vector(to_unsigned(225, 8)),
			1843 => std_logic_vector(to_unsigned(151, 8)),
			1844 => std_logic_vector(to_unsigned(66, 8)),
			1845 => std_logic_vector(to_unsigned(54, 8)),
			1846 => std_logic_vector(to_unsigned(186, 8)),
			1847 => std_logic_vector(to_unsigned(92, 8)),
			1848 => std_logic_vector(to_unsigned(30, 8)),
			1849 => std_logic_vector(to_unsigned(23, 8)),
			1850 => std_logic_vector(to_unsigned(216, 8)),
			1851 => std_logic_vector(to_unsigned(45, 8)),
			1852 => std_logic_vector(to_unsigned(198, 8)),
			1853 => std_logic_vector(to_unsigned(23, 8)),
			1854 => std_logic_vector(to_unsigned(178, 8)),
			1855 => std_logic_vector(to_unsigned(160, 8)),
			1856 => std_logic_vector(to_unsigned(141, 8)),
			1857 => std_logic_vector(to_unsigned(153, 8)),
			1858 => std_logic_vector(to_unsigned(45, 8)),
			1859 => std_logic_vector(to_unsigned(250, 8)),
			1860 => std_logic_vector(to_unsigned(29, 8)),
			1861 => std_logic_vector(to_unsigned(111, 8)),
			1862 => std_logic_vector(to_unsigned(5, 8)),
			1863 => std_logic_vector(to_unsigned(95, 8)),
			1864 => std_logic_vector(to_unsigned(205, 8)),
			1865 => std_logic_vector(to_unsigned(198, 8)),
			1866 => std_logic_vector(to_unsigned(97, 8)),
			1867 => std_logic_vector(to_unsigned(49, 8)),
			1868 => std_logic_vector(to_unsigned(137, 8)),
			1869 => std_logic_vector(to_unsigned(167, 8)),
			1870 => std_logic_vector(to_unsigned(175, 8)),
			1871 => std_logic_vector(to_unsigned(227, 8)),
			1872 => std_logic_vector(to_unsigned(252, 8)),
			1873 => std_logic_vector(to_unsigned(81, 8)),
			1874 => std_logic_vector(to_unsigned(54, 8)),
			1875 => std_logic_vector(to_unsigned(58, 8)),
			1876 => std_logic_vector(to_unsigned(63, 8)),
			1877 => std_logic_vector(to_unsigned(28, 8)),
			1878 => std_logic_vector(to_unsigned(154, 8)),
			1879 => std_logic_vector(to_unsigned(232, 8)),
			1880 => std_logic_vector(to_unsigned(133, 8)),
			1881 => std_logic_vector(to_unsigned(250, 8)),
			1882 => std_logic_vector(to_unsigned(243, 8)),
			1883 => std_logic_vector(to_unsigned(244, 8)),
			1884 => std_logic_vector(to_unsigned(29, 8)),
			1885 => std_logic_vector(to_unsigned(22, 8)),
			1886 => std_logic_vector(to_unsigned(141, 8)),
			1887 => std_logic_vector(to_unsigned(156, 8)),
			1888 => std_logic_vector(to_unsigned(107, 8)),
			1889 => std_logic_vector(to_unsigned(19, 8)),
			1890 => std_logic_vector(to_unsigned(81, 8)),
			1891 => std_logic_vector(to_unsigned(177, 8)),
			1892 => std_logic_vector(to_unsigned(166, 8)),
			1893 => std_logic_vector(to_unsigned(11, 8)),
			1894 => std_logic_vector(to_unsigned(70, 8)),
			1895 => std_logic_vector(to_unsigned(243, 8)),
			1896 => std_logic_vector(to_unsigned(239, 8)),
			1897 => std_logic_vector(to_unsigned(59, 8)),
			1898 => std_logic_vector(to_unsigned(116, 8)),
			1899 => std_logic_vector(to_unsigned(54, 8)),
			1900 => std_logic_vector(to_unsigned(99, 8)),
			1901 => std_logic_vector(to_unsigned(16, 8)),
			1902 => std_logic_vector(to_unsigned(20, 8)),
			1903 => std_logic_vector(to_unsigned(247, 8)),
			1904 => std_logic_vector(to_unsigned(199, 8)),
			1905 => std_logic_vector(to_unsigned(147, 8)),
			1906 => std_logic_vector(to_unsigned(15, 8)),
			1907 => std_logic_vector(to_unsigned(181, 8)),
			1908 => std_logic_vector(to_unsigned(120, 8)),
			1909 => std_logic_vector(to_unsigned(104, 8)),
			1910 => std_logic_vector(to_unsigned(182, 8)),
			1911 => std_logic_vector(to_unsigned(21, 8)),
			1912 => std_logic_vector(to_unsigned(231, 8)),
			1913 => std_logic_vector(to_unsigned(184, 8)),
			1914 => std_logic_vector(to_unsigned(134, 8)),
			1915 => std_logic_vector(to_unsigned(104, 8)),
			1916 => std_logic_vector(to_unsigned(21, 8)),
			1917 => std_logic_vector(to_unsigned(56, 8)),
			1918 => std_logic_vector(to_unsigned(108, 8)),
			1919 => std_logic_vector(to_unsigned(140, 8)),
			1920 => std_logic_vector(to_unsigned(4, 8)),
			1921 => std_logic_vector(to_unsigned(82, 8)),
			1922 => std_logic_vector(to_unsigned(243, 8)),
			1923 => std_logic_vector(to_unsigned(80, 8)),
			1924 => std_logic_vector(to_unsigned(163, 8)),
			1925 => std_logic_vector(to_unsigned(1, 8)),
			1926 => std_logic_vector(to_unsigned(161, 8)),
			1927 => std_logic_vector(to_unsigned(196, 8)),
			1928 => std_logic_vector(to_unsigned(129, 8)),
			1929 => std_logic_vector(to_unsigned(240, 8)),
			1930 => std_logic_vector(to_unsigned(22, 8)),
			1931 => std_logic_vector(to_unsigned(136, 8)),
			1932 => std_logic_vector(to_unsigned(141, 8)),
			1933 => std_logic_vector(to_unsigned(145, 8)),
			1934 => std_logic_vector(to_unsigned(135, 8)),
			1935 => std_logic_vector(to_unsigned(104, 8)),
			1936 => std_logic_vector(to_unsigned(129, 8)),
			1937 => std_logic_vector(to_unsigned(21, 8)),
			1938 => std_logic_vector(to_unsigned(181, 8)),
			1939 => std_logic_vector(to_unsigned(157, 8)),
			1940 => std_logic_vector(to_unsigned(194, 8)),
			1941 => std_logic_vector(to_unsigned(168, 8)),
			1942 => std_logic_vector(to_unsigned(81, 8)),
			1943 => std_logic_vector(to_unsigned(203, 8)),
			1944 => std_logic_vector(to_unsigned(241, 8)),
			1945 => std_logic_vector(to_unsigned(4, 8)),
			1946 => std_logic_vector(to_unsigned(220, 8)),
			1947 => std_logic_vector(to_unsigned(148, 8)),
			1948 => std_logic_vector(to_unsigned(210, 8)),
			1949 => std_logic_vector(to_unsigned(110, 8)),
			1950 => std_logic_vector(to_unsigned(62, 8)),
			1951 => std_logic_vector(to_unsigned(160, 8)),
			1952 => std_logic_vector(to_unsigned(227, 8)),
			1953 => std_logic_vector(to_unsigned(125, 8)),
			1954 => std_logic_vector(to_unsigned(250, 8)),
			1955 => std_logic_vector(to_unsigned(178, 8)),
			1956 => std_logic_vector(to_unsigned(136, 8)),
			1957 => std_logic_vector(to_unsigned(159, 8)),
			1958 => std_logic_vector(to_unsigned(138, 8)),
			1959 => std_logic_vector(to_unsigned(119, 8)),
			1960 => std_logic_vector(to_unsigned(236, 8)),
			1961 => std_logic_vector(to_unsigned(121, 8)),
			1962 => std_logic_vector(to_unsigned(99, 8)),
			1963 => std_logic_vector(to_unsigned(120, 8)),
			1964 => std_logic_vector(to_unsigned(12, 8)),
			1965 => std_logic_vector(to_unsigned(117, 8)),
			1966 => std_logic_vector(to_unsigned(95, 8)),
			1967 => std_logic_vector(to_unsigned(73, 8)),
			1968 => std_logic_vector(to_unsigned(160, 8)),
			1969 => std_logic_vector(to_unsigned(127, 8)),
			1970 => std_logic_vector(to_unsigned(154, 8)),
			1971 => std_logic_vector(to_unsigned(3, 8)),
			1972 => std_logic_vector(to_unsigned(196, 8)),
			1973 => std_logic_vector(to_unsigned(1, 8)),
			1974 => std_logic_vector(to_unsigned(253, 8)),
			1975 => std_logic_vector(to_unsigned(223, 8)),
			1976 => std_logic_vector(to_unsigned(40, 8)),
			1977 => std_logic_vector(to_unsigned(102, 8)),
			1978 => std_logic_vector(to_unsigned(36, 8)),
			1979 => std_logic_vector(to_unsigned(181, 8)),
			1980 => std_logic_vector(to_unsigned(0, 8)),
			1981 => std_logic_vector(to_unsigned(141, 8)),
			1982 => std_logic_vector(to_unsigned(250, 8)),
			1983 => std_logic_vector(to_unsigned(34, 8)),
			1984 => std_logic_vector(to_unsigned(240, 8)),
			1985 => std_logic_vector(to_unsigned(68, 8)),
			1986 => std_logic_vector(to_unsigned(216, 8)),
			1987 => std_logic_vector(to_unsigned(60, 8)),
			1988 => std_logic_vector(to_unsigned(50, 8)),
			1989 => std_logic_vector(to_unsigned(192, 8)),
			1990 => std_logic_vector(to_unsigned(111, 8)),
			1991 => std_logic_vector(to_unsigned(164, 8)),
			1992 => std_logic_vector(to_unsigned(54, 8)),
			1993 => std_logic_vector(to_unsigned(110, 8)),
			1994 => std_logic_vector(to_unsigned(119, 8)),
			1995 => std_logic_vector(to_unsigned(146, 8)),
			1996 => std_logic_vector(to_unsigned(91, 8)),
			1997 => std_logic_vector(to_unsigned(200, 8)),
			1998 => std_logic_vector(to_unsigned(145, 8)),
			1999 => std_logic_vector(to_unsigned(124, 8)),
			2000 => std_logic_vector(to_unsigned(193, 8)),
			2001 => std_logic_vector(to_unsigned(237, 8)),
			2002 => std_logic_vector(to_unsigned(68, 8)),
			2003 => std_logic_vector(to_unsigned(68, 8)),
			2004 => std_logic_vector(to_unsigned(47, 8)),
			2005 => std_logic_vector(to_unsigned(136, 8)),
			2006 => std_logic_vector(to_unsigned(163, 8)),
			2007 => std_logic_vector(to_unsigned(138, 8)),
			2008 => std_logic_vector(to_unsigned(42, 8)),
			2009 => std_logic_vector(to_unsigned(13, 8)),
			2010 => std_logic_vector(to_unsigned(169, 8)),
			2011 => std_logic_vector(to_unsigned(141, 8)),
			2012 => std_logic_vector(to_unsigned(211, 8)),
			2013 => std_logic_vector(to_unsigned(102, 8)),
			2014 => std_logic_vector(to_unsigned(3, 8)),
			2015 => std_logic_vector(to_unsigned(102, 8)),
			2016 => std_logic_vector(to_unsigned(58, 8)),
			2017 => std_logic_vector(to_unsigned(99, 8)),
			2018 => std_logic_vector(to_unsigned(95, 8)),
			2019 => std_logic_vector(to_unsigned(126, 8)),
			2020 => std_logic_vector(to_unsigned(77, 8)),
			2021 => std_logic_vector(to_unsigned(227, 8)),
			2022 => std_logic_vector(to_unsigned(64, 8)),
			2023 => std_logic_vector(to_unsigned(139, 8)),
			2024 => std_logic_vector(to_unsigned(230, 8)),
			2025 => std_logic_vector(to_unsigned(42, 8)),
			2026 => std_logic_vector(to_unsigned(206, 8)),
			2027 => std_logic_vector(to_unsigned(123, 8)),
			2028 => std_logic_vector(to_unsigned(131, 8)),
			2029 => std_logic_vector(to_unsigned(227, 8)),
			2030 => std_logic_vector(to_unsigned(215, 8)),
			2031 => std_logic_vector(to_unsigned(77, 8)),
			2032 => std_logic_vector(to_unsigned(8, 8)),
			2033 => std_logic_vector(to_unsigned(62, 8)),
			2034 => std_logic_vector(to_unsigned(164, 8)),
			2035 => std_logic_vector(to_unsigned(199, 8)),
			2036 => std_logic_vector(to_unsigned(66, 8)),
			2037 => std_logic_vector(to_unsigned(223, 8)),
			2038 => std_logic_vector(to_unsigned(36, 8)),
			2039 => std_logic_vector(to_unsigned(151, 8)),
			2040 => std_logic_vector(to_unsigned(100, 8)),
			2041 => std_logic_vector(to_unsigned(141, 8)),
			2042 => std_logic_vector(to_unsigned(159, 8)),
			2043 => std_logic_vector(to_unsigned(103, 8)),
			2044 => std_logic_vector(to_unsigned(131, 8)),
			2045 => std_logic_vector(to_unsigned(29, 8)),
			2046 => std_logic_vector(to_unsigned(0, 8)),
			2047 => std_logic_vector(to_unsigned(8, 8)),
			2048 => std_logic_vector(to_unsigned(254, 8)),
			2049 => std_logic_vector(to_unsigned(127, 8)),
			2050 => std_logic_vector(to_unsigned(1, 8)),
			2051 => std_logic_vector(to_unsigned(23, 8)),
			2052 => std_logic_vector(to_unsigned(165, 8)),
			2053 => std_logic_vector(to_unsigned(136, 8)),
			2054 => std_logic_vector(to_unsigned(15, 8)),
			2055 => std_logic_vector(to_unsigned(161, 8)),
			2056 => std_logic_vector(to_unsigned(161, 8)),
			2057 => std_logic_vector(to_unsigned(75, 8)),
			2058 => std_logic_vector(to_unsigned(54, 8)),
			2059 => std_logic_vector(to_unsigned(235, 8)),
			2060 => std_logic_vector(to_unsigned(143, 8)),
			2061 => std_logic_vector(to_unsigned(201, 8)),
			2062 => std_logic_vector(to_unsigned(240, 8)),
			2063 => std_logic_vector(to_unsigned(213, 8)),
			2064 => std_logic_vector(to_unsigned(133, 8)),
			2065 => std_logic_vector(to_unsigned(58, 8)),
			2066 => std_logic_vector(to_unsigned(13, 8)),
			2067 => std_logic_vector(to_unsigned(246, 8)),
			2068 => std_logic_vector(to_unsigned(49, 8)),
			2069 => std_logic_vector(to_unsigned(95, 8)),
			2070 => std_logic_vector(to_unsigned(254, 8)),
			2071 => std_logic_vector(to_unsigned(233, 8)),
			2072 => std_logic_vector(to_unsigned(220, 8)),
			2073 => std_logic_vector(to_unsigned(188, 8)),
			2074 => std_logic_vector(to_unsigned(203, 8)),
			2075 => std_logic_vector(to_unsigned(85, 8)),
			2076 => std_logic_vector(to_unsigned(101, 8)),
			2077 => std_logic_vector(to_unsigned(235, 8)),
			2078 => std_logic_vector(to_unsigned(201, 8)),
			2079 => std_logic_vector(to_unsigned(82, 8)),
			2080 => std_logic_vector(to_unsigned(141, 8)),
			2081 => std_logic_vector(to_unsigned(53, 8)),
			2082 => std_logic_vector(to_unsigned(113, 8)),
			2083 => std_logic_vector(to_unsigned(86, 8)),
			2084 => std_logic_vector(to_unsigned(221, 8)),
			2085 => std_logic_vector(to_unsigned(66, 8)),
			2086 => std_logic_vector(to_unsigned(186, 8)),
			2087 => std_logic_vector(to_unsigned(83, 8)),
			2088 => std_logic_vector(to_unsigned(15, 8)),
			2089 => std_logic_vector(to_unsigned(185, 8)),
			2090 => std_logic_vector(to_unsigned(209, 8)),
			2091 => std_logic_vector(to_unsigned(171, 8)),
			2092 => std_logic_vector(to_unsigned(191, 8)),
			2093 => std_logic_vector(to_unsigned(77, 8)),
			2094 => std_logic_vector(to_unsigned(156, 8)),
			2095 => std_logic_vector(to_unsigned(138, 8)),
			2096 => std_logic_vector(to_unsigned(88, 8)),
			2097 => std_logic_vector(to_unsigned(188, 8)),
			2098 => std_logic_vector(to_unsigned(25, 8)),
			2099 => std_logic_vector(to_unsigned(6, 8)),
			2100 => std_logic_vector(to_unsigned(220, 8)),
			2101 => std_logic_vector(to_unsigned(252, 8)),
			2102 => std_logic_vector(to_unsigned(53, 8)),
			2103 => std_logic_vector(to_unsigned(134, 8)),
			2104 => std_logic_vector(to_unsigned(84, 8)),
			2105 => std_logic_vector(to_unsigned(35, 8)),
			2106 => std_logic_vector(to_unsigned(141, 8)),
			2107 => std_logic_vector(to_unsigned(189, 8)),
			2108 => std_logic_vector(to_unsigned(99, 8)),
			2109 => std_logic_vector(to_unsigned(50, 8)),
			2110 => std_logic_vector(to_unsigned(83, 8)),
			2111 => std_logic_vector(to_unsigned(19, 8)),
			2112 => std_logic_vector(to_unsigned(176, 8)),
			2113 => std_logic_vector(to_unsigned(36, 8)),
			2114 => std_logic_vector(to_unsigned(166, 8)),
			2115 => std_logic_vector(to_unsigned(86, 8)),
			2116 => std_logic_vector(to_unsigned(6, 8)),
			2117 => std_logic_vector(to_unsigned(227, 8)),
			2118 => std_logic_vector(to_unsigned(59, 8)),
			2119 => std_logic_vector(to_unsigned(160, 8)),
			2120 => std_logic_vector(to_unsigned(84, 8)),
			2121 => std_logic_vector(to_unsigned(201, 8)),
			2122 => std_logic_vector(to_unsigned(120, 8)),
			2123 => std_logic_vector(to_unsigned(228, 8)),
			2124 => std_logic_vector(to_unsigned(232, 8)),
			2125 => std_logic_vector(to_unsigned(217, 8)),
			2126 => std_logic_vector(to_unsigned(43, 8)),
			2127 => std_logic_vector(to_unsigned(134, 8)),
			2128 => std_logic_vector(to_unsigned(33, 8)),
			2129 => std_logic_vector(to_unsigned(130, 8)),
			2130 => std_logic_vector(to_unsigned(15, 8)),
			2131 => std_logic_vector(to_unsigned(98, 8)),
			2132 => std_logic_vector(to_unsigned(82, 8)),
			2133 => std_logic_vector(to_unsigned(126, 8)),
			2134 => std_logic_vector(to_unsigned(188, 8)),
			2135 => std_logic_vector(to_unsigned(230, 8)),
			2136 => std_logic_vector(to_unsigned(253, 8)),
			2137 => std_logic_vector(to_unsigned(170, 8)),
			2138 => std_logic_vector(to_unsigned(140, 8)),
			2139 => std_logic_vector(to_unsigned(42, 8)),
			2140 => std_logic_vector(to_unsigned(157, 8)),
			2141 => std_logic_vector(to_unsigned(48, 8)),
			2142 => std_logic_vector(to_unsigned(24, 8)),
			2143 => std_logic_vector(to_unsigned(134, 8)),
			2144 => std_logic_vector(to_unsigned(103, 8)),
			2145 => std_logic_vector(to_unsigned(33, 8)),
			2146 => std_logic_vector(to_unsigned(55, 8)),
			2147 => std_logic_vector(to_unsigned(100, 8)),
			2148 => std_logic_vector(to_unsigned(242, 8)),
			2149 => std_logic_vector(to_unsigned(93, 8)),
			2150 => std_logic_vector(to_unsigned(21, 8)),
			2151 => std_logic_vector(to_unsigned(209, 8)),
			2152 => std_logic_vector(to_unsigned(254, 8)),
			2153 => std_logic_vector(to_unsigned(146, 8)),
			2154 => std_logic_vector(to_unsigned(246, 8)),
			2155 => std_logic_vector(to_unsigned(222, 8)),
			2156 => std_logic_vector(to_unsigned(201, 8)),
			2157 => std_logic_vector(to_unsigned(245, 8)),
			2158 => std_logic_vector(to_unsigned(152, 8)),
			2159 => std_logic_vector(to_unsigned(132, 8)),
			2160 => std_logic_vector(to_unsigned(42, 8)),
			2161 => std_logic_vector(to_unsigned(30, 8)),
			2162 => std_logic_vector(to_unsigned(226, 8)),
			2163 => std_logic_vector(to_unsigned(142, 8)),
			2164 => std_logic_vector(to_unsigned(229, 8)),
			2165 => std_logic_vector(to_unsigned(225, 8)),
			2166 => std_logic_vector(to_unsigned(192, 8)),
			2167 => std_logic_vector(to_unsigned(46, 8)),
			2168 => std_logic_vector(to_unsigned(91, 8)),
			2169 => std_logic_vector(to_unsigned(244, 8)),
			2170 => std_logic_vector(to_unsigned(137, 8)),
			2171 => std_logic_vector(to_unsigned(78, 8)),
			2172 => std_logic_vector(to_unsigned(159, 8)),
			2173 => std_logic_vector(to_unsigned(105, 8)),
			2174 => std_logic_vector(to_unsigned(159, 8)),
			2175 => std_logic_vector(to_unsigned(75, 8)),
			2176 => std_logic_vector(to_unsigned(27, 8)),
			2177 => std_logic_vector(to_unsigned(174, 8)),
			2178 => std_logic_vector(to_unsigned(56, 8)),
			2179 => std_logic_vector(to_unsigned(208, 8)),
			2180 => std_logic_vector(to_unsigned(45, 8)),
			2181 => std_logic_vector(to_unsigned(108, 8)),
			2182 => std_logic_vector(to_unsigned(217, 8)),
			2183 => std_logic_vector(to_unsigned(249, 8)),
			2184 => std_logic_vector(to_unsigned(211, 8)),
			2185 => std_logic_vector(to_unsigned(201, 8)),
			2186 => std_logic_vector(to_unsigned(138, 8)),
			2187 => std_logic_vector(to_unsigned(82, 8)),
			2188 => std_logic_vector(to_unsigned(213, 8)),
			2189 => std_logic_vector(to_unsigned(44, 8)),
			2190 => std_logic_vector(to_unsigned(239, 8)),
			2191 => std_logic_vector(to_unsigned(19, 8)),
			2192 => std_logic_vector(to_unsigned(198, 8)),
			2193 => std_logic_vector(to_unsigned(190, 8)),
			2194 => std_logic_vector(to_unsigned(17, 8)),
			2195 => std_logic_vector(to_unsigned(203, 8)),
			2196 => std_logic_vector(to_unsigned(99, 8)),
			2197 => std_logic_vector(to_unsigned(91, 8)),
			2198 => std_logic_vector(to_unsigned(106, 8)),
			2199 => std_logic_vector(to_unsigned(155, 8)),
			2200 => std_logic_vector(to_unsigned(186, 8)),
			2201 => std_logic_vector(to_unsigned(239, 8)),
			2202 => std_logic_vector(to_unsigned(11, 8)),
			2203 => std_logic_vector(to_unsigned(202, 8)),
			2204 => std_logic_vector(to_unsigned(194, 8)),
			2205 => std_logic_vector(to_unsigned(94, 8)),
			2206 => std_logic_vector(to_unsigned(90, 8)),
			2207 => std_logic_vector(to_unsigned(137, 8)),
			2208 => std_logic_vector(to_unsigned(8, 8)),
			2209 => std_logic_vector(to_unsigned(201, 8)),
			2210 => std_logic_vector(to_unsigned(191, 8)),
			2211 => std_logic_vector(to_unsigned(96, 8)),
			2212 => std_logic_vector(to_unsigned(201, 8)),
			2213 => std_logic_vector(to_unsigned(195, 8)),
			2214 => std_logic_vector(to_unsigned(35, 8)),
			2215 => std_logic_vector(to_unsigned(236, 8)),
			2216 => std_logic_vector(to_unsigned(100, 8)),
			2217 => std_logic_vector(to_unsigned(12, 8)),
			2218 => std_logic_vector(to_unsigned(243, 8)),
			2219 => std_logic_vector(to_unsigned(214, 8)),
			2220 => std_logic_vector(to_unsigned(163, 8)),
			2221 => std_logic_vector(to_unsigned(203, 8)),
			2222 => std_logic_vector(to_unsigned(93, 8)),
			2223 => std_logic_vector(to_unsigned(185, 8)),
			2224 => std_logic_vector(to_unsigned(36, 8)),
			2225 => std_logic_vector(to_unsigned(224, 8)),
			2226 => std_logic_vector(to_unsigned(149, 8)),
			2227 => std_logic_vector(to_unsigned(96, 8)),
			2228 => std_logic_vector(to_unsigned(133, 8)),
			2229 => std_logic_vector(to_unsigned(11, 8)),
			2230 => std_logic_vector(to_unsigned(156, 8)),
			2231 => std_logic_vector(to_unsigned(201, 8)),
			2232 => std_logic_vector(to_unsigned(60, 8)),
			2233 => std_logic_vector(to_unsigned(236, 8)),
			2234 => std_logic_vector(to_unsigned(84, 8)),
			2235 => std_logic_vector(to_unsigned(145, 8)),
			2236 => std_logic_vector(to_unsigned(255, 8)),
			2237 => std_logic_vector(to_unsigned(109, 8)),
			2238 => std_logic_vector(to_unsigned(96, 8)),
			2239 => std_logic_vector(to_unsigned(93, 8)),
			2240 => std_logic_vector(to_unsigned(94, 8)),
			2241 => std_logic_vector(to_unsigned(147, 8)),
			2242 => std_logic_vector(to_unsigned(86, 8)),
			2243 => std_logic_vector(to_unsigned(15, 8)),
			2244 => std_logic_vector(to_unsigned(20, 8)),
			2245 => std_logic_vector(to_unsigned(18, 8)),
			2246 => std_logic_vector(to_unsigned(98, 8)),
			2247 => std_logic_vector(to_unsigned(172, 8)),
			2248 => std_logic_vector(to_unsigned(173, 8)),
			2249 => std_logic_vector(to_unsigned(72, 8)),
			2250 => std_logic_vector(to_unsigned(12, 8)),
			2251 => std_logic_vector(to_unsigned(140, 8)),
			2252 => std_logic_vector(to_unsigned(195, 8)),
			2253 => std_logic_vector(to_unsigned(22, 8)),
			2254 => std_logic_vector(to_unsigned(77, 8)),
			2255 => std_logic_vector(to_unsigned(16, 8)),
			2256 => std_logic_vector(to_unsigned(143, 8)),
			2257 => std_logic_vector(to_unsigned(219, 8)),
			2258 => std_logic_vector(to_unsigned(41, 8)),
			2259 => std_logic_vector(to_unsigned(11, 8)),
			2260 => std_logic_vector(to_unsigned(187, 8)),
			2261 => std_logic_vector(to_unsigned(56, 8)),
			2262 => std_logic_vector(to_unsigned(44, 8)),
			2263 => std_logic_vector(to_unsigned(211, 8)),
			2264 => std_logic_vector(to_unsigned(205, 8)),
			2265 => std_logic_vector(to_unsigned(124, 8)),
			2266 => std_logic_vector(to_unsigned(206, 8)),
			2267 => std_logic_vector(to_unsigned(218, 8)),
			2268 => std_logic_vector(to_unsigned(94, 8)),
			2269 => std_logic_vector(to_unsigned(119, 8)),
			2270 => std_logic_vector(to_unsigned(71, 8)),
			2271 => std_logic_vector(to_unsigned(44, 8)),
			2272 => std_logic_vector(to_unsigned(227, 8)),
			2273 => std_logic_vector(to_unsigned(135, 8)),
			2274 => std_logic_vector(to_unsigned(220, 8)),
			2275 => std_logic_vector(to_unsigned(62, 8)),
			2276 => std_logic_vector(to_unsigned(216, 8)),
			2277 => std_logic_vector(to_unsigned(134, 8)),
			2278 => std_logic_vector(to_unsigned(183, 8)),
			2279 => std_logic_vector(to_unsigned(28, 8)),
			2280 => std_logic_vector(to_unsigned(7, 8)),
			2281 => std_logic_vector(to_unsigned(28, 8)),
			2282 => std_logic_vector(to_unsigned(175, 8)),
			2283 => std_logic_vector(to_unsigned(248, 8)),
			2284 => std_logic_vector(to_unsigned(79, 8)),
			2285 => std_logic_vector(to_unsigned(138, 8)),
			2286 => std_logic_vector(to_unsigned(55, 8)),
			2287 => std_logic_vector(to_unsigned(234, 8)),
			2288 => std_logic_vector(to_unsigned(61, 8)),
			2289 => std_logic_vector(to_unsigned(31, 8)),
			2290 => std_logic_vector(to_unsigned(165, 8)),
			2291 => std_logic_vector(to_unsigned(43, 8)),
			2292 => std_logic_vector(to_unsigned(175, 8)),
			2293 => std_logic_vector(to_unsigned(231, 8)),
			2294 => std_logic_vector(to_unsigned(222, 8)),
			2295 => std_logic_vector(to_unsigned(222, 8)),
			2296 => std_logic_vector(to_unsigned(101, 8)),
			2297 => std_logic_vector(to_unsigned(190, 8)),
			2298 => std_logic_vector(to_unsigned(240, 8)),
			2299 => std_logic_vector(to_unsigned(89, 8)),
			2300 => std_logic_vector(to_unsigned(3, 8)),
			2301 => std_logic_vector(to_unsigned(102, 8)),
			2302 => std_logic_vector(to_unsigned(143, 8)),
			2303 => std_logic_vector(to_unsigned(27, 8)),
			2304 => std_logic_vector(to_unsigned(5, 8)),
			2305 => std_logic_vector(to_unsigned(100, 8)),
			2306 => std_logic_vector(to_unsigned(79, 8)),
			2307 => std_logic_vector(to_unsigned(73, 8)),
			2308 => std_logic_vector(to_unsigned(103, 8)),
			2309 => std_logic_vector(to_unsigned(129, 8)),
			2310 => std_logic_vector(to_unsigned(88, 8)),
			2311 => std_logic_vector(to_unsigned(72, 8)),
			2312 => std_logic_vector(to_unsigned(160, 8)),
			2313 => std_logic_vector(to_unsigned(237, 8)),
			2314 => std_logic_vector(to_unsigned(37, 8)),
			2315 => std_logic_vector(to_unsigned(93, 8)),
			2316 => std_logic_vector(to_unsigned(217, 8)),
			2317 => std_logic_vector(to_unsigned(214, 8)),
			2318 => std_logic_vector(to_unsigned(73, 8)),
			2319 => std_logic_vector(to_unsigned(196, 8)),
			2320 => std_logic_vector(to_unsigned(20, 8)),
			2321 => std_logic_vector(to_unsigned(226, 8)),
			2322 => std_logic_vector(to_unsigned(218, 8)),
			2323 => std_logic_vector(to_unsigned(164, 8)),
			2324 => std_logic_vector(to_unsigned(172, 8)),
			2325 => std_logic_vector(to_unsigned(20, 8)),
			2326 => std_logic_vector(to_unsigned(176, 8)),
			2327 => std_logic_vector(to_unsigned(206, 8)),
			2328 => std_logic_vector(to_unsigned(68, 8)),
			2329 => std_logic_vector(to_unsigned(253, 8)),
			2330 => std_logic_vector(to_unsigned(160, 8)),
			2331 => std_logic_vector(to_unsigned(179, 8)),
			2332 => std_logic_vector(to_unsigned(102, 8)),
			2333 => std_logic_vector(to_unsigned(48, 8)),
			2334 => std_logic_vector(to_unsigned(8, 8)),
			2335 => std_logic_vector(to_unsigned(141, 8)),
			2336 => std_logic_vector(to_unsigned(243, 8)),
			2337 => std_logic_vector(to_unsigned(173, 8)),
			2338 => std_logic_vector(to_unsigned(56, 8)),
			2339 => std_logic_vector(to_unsigned(220, 8)),
			2340 => std_logic_vector(to_unsigned(235, 8)),
			2341 => std_logic_vector(to_unsigned(101, 8)),
			2342 => std_logic_vector(to_unsigned(8, 8)),
			2343 => std_logic_vector(to_unsigned(132, 8)),
			2344 => std_logic_vector(to_unsigned(32, 8)),
			2345 => std_logic_vector(to_unsigned(84, 8)),
			2346 => std_logic_vector(to_unsigned(185, 8)),
			2347 => std_logic_vector(to_unsigned(113, 8)),
			2348 => std_logic_vector(to_unsigned(5, 8)),
			2349 => std_logic_vector(to_unsigned(247, 8)),
			2350 => std_logic_vector(to_unsigned(94, 8)),
			2351 => std_logic_vector(to_unsigned(178, 8)),
			2352 => std_logic_vector(to_unsigned(206, 8)),
			2353 => std_logic_vector(to_unsigned(146, 8)),
			2354 => std_logic_vector(to_unsigned(128, 8)),
			2355 => std_logic_vector(to_unsigned(101, 8)),
			2356 => std_logic_vector(to_unsigned(210, 8)),
			2357 => std_logic_vector(to_unsigned(212, 8)),
			2358 => std_logic_vector(to_unsigned(228, 8)),
			2359 => std_logic_vector(to_unsigned(74, 8)),
			2360 => std_logic_vector(to_unsigned(199, 8)),
			2361 => std_logic_vector(to_unsigned(144, 8)),
			2362 => std_logic_vector(to_unsigned(14, 8)),
			2363 => std_logic_vector(to_unsigned(70, 8)),
			2364 => std_logic_vector(to_unsigned(179, 8)),
			2365 => std_logic_vector(to_unsigned(169, 8)),
			2366 => std_logic_vector(to_unsigned(181, 8)),
			2367 => std_logic_vector(to_unsigned(171, 8)),
			2368 => std_logic_vector(to_unsigned(147, 8)),
			2369 => std_logic_vector(to_unsigned(170, 8)),
			2370 => std_logic_vector(to_unsigned(242, 8)),
			2371 => std_logic_vector(to_unsigned(41, 8)),
			2372 => std_logic_vector(to_unsigned(202, 8)),
			2373 => std_logic_vector(to_unsigned(25, 8)),
			2374 => std_logic_vector(to_unsigned(198, 8)),
			2375 => std_logic_vector(to_unsigned(120, 8)),
			2376 => std_logic_vector(to_unsigned(90, 8)),
			2377 => std_logic_vector(to_unsigned(56, 8)),
			2378 => std_logic_vector(to_unsigned(24, 8)),
			2379 => std_logic_vector(to_unsigned(123, 8)),
			2380 => std_logic_vector(to_unsigned(92, 8)),
			2381 => std_logic_vector(to_unsigned(52, 8)),
			2382 => std_logic_vector(to_unsigned(132, 8)),
			2383 => std_logic_vector(to_unsigned(102, 8)),
			2384 => std_logic_vector(to_unsigned(129, 8)),
			2385 => std_logic_vector(to_unsigned(121, 8)),
			2386 => std_logic_vector(to_unsigned(254, 8)),
			2387 => std_logic_vector(to_unsigned(188, 8)),
			2388 => std_logic_vector(to_unsigned(218, 8)),
			2389 => std_logic_vector(to_unsigned(18, 8)),
			2390 => std_logic_vector(to_unsigned(250, 8)),
			2391 => std_logic_vector(to_unsigned(0, 8)),
			2392 => std_logic_vector(to_unsigned(32, 8)),
			2393 => std_logic_vector(to_unsigned(166, 8)),
			2394 => std_logic_vector(to_unsigned(240, 8)),
			2395 => std_logic_vector(to_unsigned(35, 8)),
			2396 => std_logic_vector(to_unsigned(50, 8)),
			2397 => std_logic_vector(to_unsigned(19, 8)),
			2398 => std_logic_vector(to_unsigned(43, 8)),
			2399 => std_logic_vector(to_unsigned(169, 8)),
			2400 => std_logic_vector(to_unsigned(152, 8)),
			2401 => std_logic_vector(to_unsigned(26, 8)),
			2402 => std_logic_vector(to_unsigned(247, 8)),
			2403 => std_logic_vector(to_unsigned(215, 8)),
			2404 => std_logic_vector(to_unsigned(35, 8)),
			2405 => std_logic_vector(to_unsigned(175, 8)),
			2406 => std_logic_vector(to_unsigned(82, 8)),
			2407 => std_logic_vector(to_unsigned(210, 8)),
			2408 => std_logic_vector(to_unsigned(173, 8)),
			2409 => std_logic_vector(to_unsigned(150, 8)),
			2410 => std_logic_vector(to_unsigned(108, 8)),
			2411 => std_logic_vector(to_unsigned(163, 8)),
			2412 => std_logic_vector(to_unsigned(217, 8)),
			2413 => std_logic_vector(to_unsigned(54, 8)),
			2414 => std_logic_vector(to_unsigned(147, 8)),
			2415 => std_logic_vector(to_unsigned(212, 8)),
			2416 => std_logic_vector(to_unsigned(61, 8)),
			2417 => std_logic_vector(to_unsigned(220, 8)),
			2418 => std_logic_vector(to_unsigned(138, 8)),
			2419 => std_logic_vector(to_unsigned(95, 8)),
			2420 => std_logic_vector(to_unsigned(103, 8)),
			2421 => std_logic_vector(to_unsigned(56, 8)),
			2422 => std_logic_vector(to_unsigned(147, 8)),
			2423 => std_logic_vector(to_unsigned(237, 8)),
			2424 => std_logic_vector(to_unsigned(109, 8)),
			2425 => std_logic_vector(to_unsigned(56, 8)),
			2426 => std_logic_vector(to_unsigned(51, 8)),
			2427 => std_logic_vector(to_unsigned(101, 8)),
			2428 => std_logic_vector(to_unsigned(83, 8)),
			2429 => std_logic_vector(to_unsigned(80, 8)),
			2430 => std_logic_vector(to_unsigned(191, 8)),
			2431 => std_logic_vector(to_unsigned(188, 8)),
			2432 => std_logic_vector(to_unsigned(171, 8)),
			2433 => std_logic_vector(to_unsigned(220, 8)),
			2434 => std_logic_vector(to_unsigned(132, 8)),
			2435 => std_logic_vector(to_unsigned(228, 8)),
			2436 => std_logic_vector(to_unsigned(32, 8)),
			2437 => std_logic_vector(to_unsigned(51, 8)),
			2438 => std_logic_vector(to_unsigned(83, 8)),
			2439 => std_logic_vector(to_unsigned(90, 8)),
			2440 => std_logic_vector(to_unsigned(62, 8)),
			2441 => std_logic_vector(to_unsigned(131, 8)),
			2442 => std_logic_vector(to_unsigned(239, 8)),
			2443 => std_logic_vector(to_unsigned(44, 8)),
			2444 => std_logic_vector(to_unsigned(125, 8)),
			2445 => std_logic_vector(to_unsigned(69, 8)),
			2446 => std_logic_vector(to_unsigned(24, 8)),
			2447 => std_logic_vector(to_unsigned(220, 8)),
			2448 => std_logic_vector(to_unsigned(115, 8)),
			2449 => std_logic_vector(to_unsigned(237, 8)),
			2450 => std_logic_vector(to_unsigned(128, 8)),
			2451 => std_logic_vector(to_unsigned(156, 8)),
			2452 => std_logic_vector(to_unsigned(120, 8)),
			2453 => std_logic_vector(to_unsigned(249, 8)),
			2454 => std_logic_vector(to_unsigned(184, 8)),
			2455 => std_logic_vector(to_unsigned(191, 8)),
			2456 => std_logic_vector(to_unsigned(73, 8)),
			2457 => std_logic_vector(to_unsigned(254, 8)),
			2458 => std_logic_vector(to_unsigned(141, 8)),
			2459 => std_logic_vector(to_unsigned(203, 8)),
			2460 => std_logic_vector(to_unsigned(124, 8)),
			2461 => std_logic_vector(to_unsigned(231, 8)),
			2462 => std_logic_vector(to_unsigned(148, 8)),
			2463 => std_logic_vector(to_unsigned(96, 8)),
			2464 => std_logic_vector(to_unsigned(203, 8)),
			2465 => std_logic_vector(to_unsigned(76, 8)),
			2466 => std_logic_vector(to_unsigned(183, 8)),
			2467 => std_logic_vector(to_unsigned(83, 8)),
			2468 => std_logic_vector(to_unsigned(47, 8)),
			2469 => std_logic_vector(to_unsigned(98, 8)),
			2470 => std_logic_vector(to_unsigned(57, 8)),
			2471 => std_logic_vector(to_unsigned(177, 8)),
			2472 => std_logic_vector(to_unsigned(176, 8)),
			2473 => std_logic_vector(to_unsigned(16, 8)),
			2474 => std_logic_vector(to_unsigned(117, 8)),
			2475 => std_logic_vector(to_unsigned(112, 8)),
			2476 => std_logic_vector(to_unsigned(247, 8)),
			2477 => std_logic_vector(to_unsigned(48, 8)),
			2478 => std_logic_vector(to_unsigned(30, 8)),
			2479 => std_logic_vector(to_unsigned(157, 8)),
			2480 => std_logic_vector(to_unsigned(131, 8)),
			2481 => std_logic_vector(to_unsigned(49, 8)),
			2482 => std_logic_vector(to_unsigned(235, 8)),
			2483 => std_logic_vector(to_unsigned(158, 8)),
			2484 => std_logic_vector(to_unsigned(33, 8)),
			2485 => std_logic_vector(to_unsigned(107, 8)),
			2486 => std_logic_vector(to_unsigned(254, 8)),
			2487 => std_logic_vector(to_unsigned(217, 8)),
			2488 => std_logic_vector(to_unsigned(198, 8)),
			2489 => std_logic_vector(to_unsigned(204, 8)),
			2490 => std_logic_vector(to_unsigned(81, 8)),
			2491 => std_logic_vector(to_unsigned(44, 8)),
			2492 => std_logic_vector(to_unsigned(207, 8)),
			2493 => std_logic_vector(to_unsigned(101, 8)),
			2494 => std_logic_vector(to_unsigned(233, 8)),
			2495 => std_logic_vector(to_unsigned(8, 8)),
			2496 => std_logic_vector(to_unsigned(251, 8)),
			2497 => std_logic_vector(to_unsigned(251, 8)),
			2498 => std_logic_vector(to_unsigned(4, 8)),
			2499 => std_logic_vector(to_unsigned(73, 8)),
			2500 => std_logic_vector(to_unsigned(82, 8)),
			2501 => std_logic_vector(to_unsigned(237, 8)),
			2502 => std_logic_vector(to_unsigned(140, 8)),
			2503 => std_logic_vector(to_unsigned(152, 8)),
			2504 => std_logic_vector(to_unsigned(218, 8)),
			2505 => std_logic_vector(to_unsigned(184, 8)),
			2506 => std_logic_vector(to_unsigned(76, 8)),
			2507 => std_logic_vector(to_unsigned(90, 8)),
			2508 => std_logic_vector(to_unsigned(176, 8)),
			2509 => std_logic_vector(to_unsigned(217, 8)),
			2510 => std_logic_vector(to_unsigned(218, 8)),
			2511 => std_logic_vector(to_unsigned(254, 8)),
			2512 => std_logic_vector(to_unsigned(69, 8)),
			2513 => std_logic_vector(to_unsigned(244, 8)),
			2514 => std_logic_vector(to_unsigned(161, 8)),
			2515 => std_logic_vector(to_unsigned(153, 8)),
			2516 => std_logic_vector(to_unsigned(156, 8)),
			2517 => std_logic_vector(to_unsigned(197, 8)),
			2518 => std_logic_vector(to_unsigned(190, 8)),
			2519 => std_logic_vector(to_unsigned(242, 8)),
			2520 => std_logic_vector(to_unsigned(222, 8)),
			2521 => std_logic_vector(to_unsigned(227, 8)),
			2522 => std_logic_vector(to_unsigned(197, 8)),
			2523 => std_logic_vector(to_unsigned(157, 8)),
			2524 => std_logic_vector(to_unsigned(22, 8)),
			2525 => std_logic_vector(to_unsigned(19, 8)),
			2526 => std_logic_vector(to_unsigned(254, 8)),
			2527 => std_logic_vector(to_unsigned(110, 8)),
			2528 => std_logic_vector(to_unsigned(113, 8)),
			2529 => std_logic_vector(to_unsigned(159, 8)),
			2530 => std_logic_vector(to_unsigned(138, 8)),
			2531 => std_logic_vector(to_unsigned(166, 8)),
			2532 => std_logic_vector(to_unsigned(10, 8)),
			2533 => std_logic_vector(to_unsigned(187, 8)),
			2534 => std_logic_vector(to_unsigned(71, 8)),
			2535 => std_logic_vector(to_unsigned(172, 8)),
			2536 => std_logic_vector(to_unsigned(178, 8)),
			2537 => std_logic_vector(to_unsigned(38, 8)),
			2538 => std_logic_vector(to_unsigned(188, 8)),
			2539 => std_logic_vector(to_unsigned(142, 8)),
			2540 => std_logic_vector(to_unsigned(98, 8)),
			2541 => std_logic_vector(to_unsigned(39, 8)),
			2542 => std_logic_vector(to_unsigned(78, 8)),
			2543 => std_logic_vector(to_unsigned(117, 8)),
			2544 => std_logic_vector(to_unsigned(247, 8)),
			2545 => std_logic_vector(to_unsigned(58, 8)),
			2546 => std_logic_vector(to_unsigned(210, 8)),
			2547 => std_logic_vector(to_unsigned(2, 8)),
			2548 => std_logic_vector(to_unsigned(84, 8)),
			2549 => std_logic_vector(to_unsigned(120, 8)),
			2550 => std_logic_vector(to_unsigned(8, 8)),
			2551 => std_logic_vector(to_unsigned(180, 8)),
			2552 => std_logic_vector(to_unsigned(252, 8)),
			2553 => std_logic_vector(to_unsigned(39, 8)),
			2554 => std_logic_vector(to_unsigned(116, 8)),
			2555 => std_logic_vector(to_unsigned(120, 8)),
			2556 => std_logic_vector(to_unsigned(143, 8)),
			2557 => std_logic_vector(to_unsigned(64, 8)),
			2558 => std_logic_vector(to_unsigned(149, 8)),
			2559 => std_logic_vector(to_unsigned(21, 8)),
			2560 => std_logic_vector(to_unsigned(138, 8)),
			2561 => std_logic_vector(to_unsigned(5, 8)),
			2562 => std_logic_vector(to_unsigned(137, 8)),
			2563 => std_logic_vector(to_unsigned(201, 8)),
			2564 => std_logic_vector(to_unsigned(171, 8)),
			2565 => std_logic_vector(to_unsigned(133, 8)),
			2566 => std_logic_vector(to_unsigned(133, 8)),
			2567 => std_logic_vector(to_unsigned(173, 8)),
			2568 => std_logic_vector(to_unsigned(52, 8)),
			2569 => std_logic_vector(to_unsigned(7, 8)),
			2570 => std_logic_vector(to_unsigned(112, 8)),
			2571 => std_logic_vector(to_unsigned(129, 8)),
			2572 => std_logic_vector(to_unsigned(137, 8)),
			2573 => std_logic_vector(to_unsigned(154, 8)),
			2574 => std_logic_vector(to_unsigned(77, 8)),
			2575 => std_logic_vector(to_unsigned(151, 8)),
			2576 => std_logic_vector(to_unsigned(255, 8)),
			2577 => std_logic_vector(to_unsigned(185, 8)),
			2578 => std_logic_vector(to_unsigned(43, 8)),
			2579 => std_logic_vector(to_unsigned(226, 8)),
			2580 => std_logic_vector(to_unsigned(221, 8)),
			2581 => std_logic_vector(to_unsigned(21, 8)),
			2582 => std_logic_vector(to_unsigned(220, 8)),
			2583 => std_logic_vector(to_unsigned(55, 8)),
			2584 => std_logic_vector(to_unsigned(12, 8)),
			2585 => std_logic_vector(to_unsigned(144, 8)),
			2586 => std_logic_vector(to_unsigned(213, 8)),
			2587 => std_logic_vector(to_unsigned(73, 8)),
			2588 => std_logic_vector(to_unsigned(156, 8)),
			2589 => std_logic_vector(to_unsigned(90, 8)),
			2590 => std_logic_vector(to_unsigned(15, 8)),
			2591 => std_logic_vector(to_unsigned(154, 8)),
			2592 => std_logic_vector(to_unsigned(44, 8)),
			2593 => std_logic_vector(to_unsigned(130, 8)),
			2594 => std_logic_vector(to_unsigned(136, 8)),
			2595 => std_logic_vector(to_unsigned(215, 8)),
			2596 => std_logic_vector(to_unsigned(85, 8)),
			2597 => std_logic_vector(to_unsigned(161, 8)),
			2598 => std_logic_vector(to_unsigned(53, 8)),
			2599 => std_logic_vector(to_unsigned(168, 8)),
			2600 => std_logic_vector(to_unsigned(22, 8)),
			2601 => std_logic_vector(to_unsigned(246, 8)),
			2602 => std_logic_vector(to_unsigned(189, 8)),
			2603 => std_logic_vector(to_unsigned(216, 8)),
			2604 => std_logic_vector(to_unsigned(241, 8)),
			2605 => std_logic_vector(to_unsigned(203, 8)),
			2606 => std_logic_vector(to_unsigned(251, 8)),
			2607 => std_logic_vector(to_unsigned(86, 8)),
			2608 => std_logic_vector(to_unsigned(206, 8)),
			2609 => std_logic_vector(to_unsigned(142, 8)),
			2610 => std_logic_vector(to_unsigned(121, 8)),
			2611 => std_logic_vector(to_unsigned(192, 8)),
			2612 => std_logic_vector(to_unsigned(30, 8)),
			2613 => std_logic_vector(to_unsigned(87, 8)),
			2614 => std_logic_vector(to_unsigned(108, 8)),
			2615 => std_logic_vector(to_unsigned(117, 8)),
			2616 => std_logic_vector(to_unsigned(147, 8)),
			2617 => std_logic_vector(to_unsigned(96, 8)),
			2618 => std_logic_vector(to_unsigned(164, 8)),
			2619 => std_logic_vector(to_unsigned(248, 8)),
			2620 => std_logic_vector(to_unsigned(227, 8)),
			2621 => std_logic_vector(to_unsigned(228, 8)),
			2622 => std_logic_vector(to_unsigned(93, 8)),
			2623 => std_logic_vector(to_unsigned(172, 8)),
			2624 => std_logic_vector(to_unsigned(236, 8)),
			2625 => std_logic_vector(to_unsigned(174, 8)),
			2626 => std_logic_vector(to_unsigned(34, 8)),
			2627 => std_logic_vector(to_unsigned(106, 8)),
			2628 => std_logic_vector(to_unsigned(70, 8)),
			2629 => std_logic_vector(to_unsigned(43, 8)),
			2630 => std_logic_vector(to_unsigned(150, 8)),
			2631 => std_logic_vector(to_unsigned(180, 8)),
			2632 => std_logic_vector(to_unsigned(133, 8)),
			2633 => std_logic_vector(to_unsigned(215, 8)),
			2634 => std_logic_vector(to_unsigned(53, 8)),
			2635 => std_logic_vector(to_unsigned(45, 8)),
			2636 => std_logic_vector(to_unsigned(14, 8)),
			2637 => std_logic_vector(to_unsigned(111, 8)),
			2638 => std_logic_vector(to_unsigned(235, 8)),
			2639 => std_logic_vector(to_unsigned(156, 8)),
			2640 => std_logic_vector(to_unsigned(177, 8)),
			2641 => std_logic_vector(to_unsigned(235, 8)),
			2642 => std_logic_vector(to_unsigned(137, 8)),
			2643 => std_logic_vector(to_unsigned(193, 8)),
			2644 => std_logic_vector(to_unsigned(42, 8)),
			2645 => std_logic_vector(to_unsigned(12, 8)),
			2646 => std_logic_vector(to_unsigned(6, 8)),
			2647 => std_logic_vector(to_unsigned(229, 8)),
			2648 => std_logic_vector(to_unsigned(14, 8)),
			2649 => std_logic_vector(to_unsigned(124, 8)),
			2650 => std_logic_vector(to_unsigned(182, 8)),
			2651 => std_logic_vector(to_unsigned(42, 8)),
			2652 => std_logic_vector(to_unsigned(105, 8)),
			2653 => std_logic_vector(to_unsigned(42, 8)),
			2654 => std_logic_vector(to_unsigned(121, 8)),
			2655 => std_logic_vector(to_unsigned(158, 8)),
			2656 => std_logic_vector(to_unsigned(130, 8)),
			2657 => std_logic_vector(to_unsigned(32, 8)),
			2658 => std_logic_vector(to_unsigned(194, 8)),
			2659 => std_logic_vector(to_unsigned(89, 8)),
			2660 => std_logic_vector(to_unsigned(86, 8)),
			2661 => std_logic_vector(to_unsigned(52, 8)),
			2662 => std_logic_vector(to_unsigned(49, 8)),
			2663 => std_logic_vector(to_unsigned(180, 8)),
			2664 => std_logic_vector(to_unsigned(114, 8)),
			2665 => std_logic_vector(to_unsigned(178, 8)),
			2666 => std_logic_vector(to_unsigned(166, 8)),
			2667 => std_logic_vector(to_unsigned(197, 8)),
			2668 => std_logic_vector(to_unsigned(209, 8)),
			2669 => std_logic_vector(to_unsigned(84, 8)),
			2670 => std_logic_vector(to_unsigned(60, 8)),
			2671 => std_logic_vector(to_unsigned(198, 8)),
			2672 => std_logic_vector(to_unsigned(235, 8)),
			2673 => std_logic_vector(to_unsigned(122, 8)),
			2674 => std_logic_vector(to_unsigned(78, 8)),
			2675 => std_logic_vector(to_unsigned(251, 8)),
			2676 => std_logic_vector(to_unsigned(2, 8)),
			2677 => std_logic_vector(to_unsigned(80, 8)),
			2678 => std_logic_vector(to_unsigned(230, 8)),
			2679 => std_logic_vector(to_unsigned(196, 8)),
			2680 => std_logic_vector(to_unsigned(156, 8)),
			2681 => std_logic_vector(to_unsigned(203, 8)),
			2682 => std_logic_vector(to_unsigned(25, 8)),
			2683 => std_logic_vector(to_unsigned(224, 8)),
			2684 => std_logic_vector(to_unsigned(175, 8)),
			2685 => std_logic_vector(to_unsigned(121, 8)),
			2686 => std_logic_vector(to_unsigned(181, 8)),
			2687 => std_logic_vector(to_unsigned(54, 8)),
			2688 => std_logic_vector(to_unsigned(205, 8)),
			2689 => std_logic_vector(to_unsigned(108, 8)),
			2690 => std_logic_vector(to_unsigned(255, 8)),
			2691 => std_logic_vector(to_unsigned(123, 8)),
			2692 => std_logic_vector(to_unsigned(78, 8)),
			2693 => std_logic_vector(to_unsigned(36, 8)),
			2694 => std_logic_vector(to_unsigned(167, 8)),
			2695 => std_logic_vector(to_unsigned(15, 8)),
			2696 => std_logic_vector(to_unsigned(74, 8)),
			2697 => std_logic_vector(to_unsigned(102, 8)),
			2698 => std_logic_vector(to_unsigned(169, 8)),
			2699 => std_logic_vector(to_unsigned(29, 8)),
			2700 => std_logic_vector(to_unsigned(64, 8)),
			2701 => std_logic_vector(to_unsigned(121, 8)),
			2702 => std_logic_vector(to_unsigned(187, 8)),
			2703 => std_logic_vector(to_unsigned(17, 8)),
			2704 => std_logic_vector(to_unsigned(116, 8)),
			2705 => std_logic_vector(to_unsigned(254, 8)),
			2706 => std_logic_vector(to_unsigned(174, 8)),
			2707 => std_logic_vector(to_unsigned(118, 8)),
			2708 => std_logic_vector(to_unsigned(238, 8)),
			2709 => std_logic_vector(to_unsigned(64, 8)),
			2710 => std_logic_vector(to_unsigned(57, 8)),
			2711 => std_logic_vector(to_unsigned(72, 8)),
			2712 => std_logic_vector(to_unsigned(66, 8)),
			2713 => std_logic_vector(to_unsigned(229, 8)),
			2714 => std_logic_vector(to_unsigned(47, 8)),
			2715 => std_logic_vector(to_unsigned(209, 8)),
			2716 => std_logic_vector(to_unsigned(69, 8)),
			2717 => std_logic_vector(to_unsigned(91, 8)),
			2718 => std_logic_vector(to_unsigned(232, 8)),
			2719 => std_logic_vector(to_unsigned(107, 8)),
			2720 => std_logic_vector(to_unsigned(244, 8)),
			2721 => std_logic_vector(to_unsigned(14, 8)),
			2722 => std_logic_vector(to_unsigned(47, 8)),
			2723 => std_logic_vector(to_unsigned(169, 8)),
			2724 => std_logic_vector(to_unsigned(101, 8)),
			2725 => std_logic_vector(to_unsigned(171, 8)),
			2726 => std_logic_vector(to_unsigned(218, 8)),
			2727 => std_logic_vector(to_unsigned(26, 8)),
			2728 => std_logic_vector(to_unsigned(180, 8)),
			2729 => std_logic_vector(to_unsigned(62, 8)),
			2730 => std_logic_vector(to_unsigned(251, 8)),
			2731 => std_logic_vector(to_unsigned(150, 8)),
			2732 => std_logic_vector(to_unsigned(163, 8)),
			2733 => std_logic_vector(to_unsigned(66, 8)),
			2734 => std_logic_vector(to_unsigned(194, 8)),
			2735 => std_logic_vector(to_unsigned(137, 8)),
			2736 => std_logic_vector(to_unsigned(186, 8)),
			2737 => std_logic_vector(to_unsigned(96, 8)),
			2738 => std_logic_vector(to_unsigned(100, 8)),
			2739 => std_logic_vector(to_unsigned(65, 8)),
			2740 => std_logic_vector(to_unsigned(36, 8)),
			2741 => std_logic_vector(to_unsigned(95, 8)),
			2742 => std_logic_vector(to_unsigned(36, 8)),
			2743 => std_logic_vector(to_unsigned(63, 8)),
			2744 => std_logic_vector(to_unsigned(47, 8)),
			2745 => std_logic_vector(to_unsigned(174, 8)),
			2746 => std_logic_vector(to_unsigned(208, 8)),
			2747 => std_logic_vector(to_unsigned(185, 8)),
			2748 => std_logic_vector(to_unsigned(199, 8)),
			2749 => std_logic_vector(to_unsigned(157, 8)),
			2750 => std_logic_vector(to_unsigned(1, 8)),
			2751 => std_logic_vector(to_unsigned(188, 8)),
			2752 => std_logic_vector(to_unsigned(168, 8)),
			2753 => std_logic_vector(to_unsigned(245, 8)),
			2754 => std_logic_vector(to_unsigned(42, 8)),
			2755 => std_logic_vector(to_unsigned(146, 8)),
			2756 => std_logic_vector(to_unsigned(83, 8)),
			2757 => std_logic_vector(to_unsigned(159, 8)),
			2758 => std_logic_vector(to_unsigned(187, 8)),
			2759 => std_logic_vector(to_unsigned(58, 8)),
			2760 => std_logic_vector(to_unsigned(92, 8)),
			2761 => std_logic_vector(to_unsigned(30, 8)),
			2762 => std_logic_vector(to_unsigned(115, 8)),
			2763 => std_logic_vector(to_unsigned(195, 8)),
			2764 => std_logic_vector(to_unsigned(106, 8)),
			2765 => std_logic_vector(to_unsigned(248, 8)),
			2766 => std_logic_vector(to_unsigned(103, 8)),
			2767 => std_logic_vector(to_unsigned(204, 8)),
			2768 => std_logic_vector(to_unsigned(139, 8)),
			2769 => std_logic_vector(to_unsigned(49, 8)),
			2770 => std_logic_vector(to_unsigned(37, 8)),
			2771 => std_logic_vector(to_unsigned(23, 8)),
			2772 => std_logic_vector(to_unsigned(162, 8)),
			2773 => std_logic_vector(to_unsigned(222, 8)),
			2774 => std_logic_vector(to_unsigned(210, 8)),
			2775 => std_logic_vector(to_unsigned(131, 8)),
			2776 => std_logic_vector(to_unsigned(197, 8)),
			2777 => std_logic_vector(to_unsigned(208, 8)),
			2778 => std_logic_vector(to_unsigned(143, 8)),
			2779 => std_logic_vector(to_unsigned(149, 8)),
			2780 => std_logic_vector(to_unsigned(59, 8)),
			2781 => std_logic_vector(to_unsigned(160, 8)),
			2782 => std_logic_vector(to_unsigned(125, 8)),
			2783 => std_logic_vector(to_unsigned(140, 8)),
			2784 => std_logic_vector(to_unsigned(164, 8)),
			2785 => std_logic_vector(to_unsigned(118, 8)),
			2786 => std_logic_vector(to_unsigned(127, 8)),
			2787 => std_logic_vector(to_unsigned(162, 8)),
			2788 => std_logic_vector(to_unsigned(140, 8)),
			2789 => std_logic_vector(to_unsigned(70, 8)),
			2790 => std_logic_vector(to_unsigned(217, 8)),
			2791 => std_logic_vector(to_unsigned(143, 8)),
			2792 => std_logic_vector(to_unsigned(159, 8)),
			2793 => std_logic_vector(to_unsigned(224, 8)),
			2794 => std_logic_vector(to_unsigned(134, 8)),
			2795 => std_logic_vector(to_unsigned(124, 8)),
			2796 => std_logic_vector(to_unsigned(77, 8)),
			2797 => std_logic_vector(to_unsigned(72, 8)),
			2798 => std_logic_vector(to_unsigned(13, 8)),
			2799 => std_logic_vector(to_unsigned(58, 8)),
			2800 => std_logic_vector(to_unsigned(52, 8)),
			2801 => std_logic_vector(to_unsigned(110, 8)),
			2802 => std_logic_vector(to_unsigned(78, 8)),
			2803 => std_logic_vector(to_unsigned(186, 8)),
			2804 => std_logic_vector(to_unsigned(171, 8)),
			2805 => std_logic_vector(to_unsigned(249, 8)),
			2806 => std_logic_vector(to_unsigned(201, 8)),
			2807 => std_logic_vector(to_unsigned(30, 8)),
			2808 => std_logic_vector(to_unsigned(180, 8)),
			2809 => std_logic_vector(to_unsigned(197, 8)),
			2810 => std_logic_vector(to_unsigned(200, 8)),
			2811 => std_logic_vector(to_unsigned(202, 8)),
			2812 => std_logic_vector(to_unsigned(136, 8)),
			2813 => std_logic_vector(to_unsigned(177, 8)),
			2814 => std_logic_vector(to_unsigned(204, 8)),
			2815 => std_logic_vector(to_unsigned(135, 8)),
			2816 => std_logic_vector(to_unsigned(237, 8)),
			2817 => std_logic_vector(to_unsigned(176, 8)),
			2818 => std_logic_vector(to_unsigned(12, 8)),
			2819 => std_logic_vector(to_unsigned(198, 8)),
			2820 => std_logic_vector(to_unsigned(25, 8)),
			2821 => std_logic_vector(to_unsigned(54, 8)),
			2822 => std_logic_vector(to_unsigned(201, 8)),
			2823 => std_logic_vector(to_unsigned(23, 8)),
			2824 => std_logic_vector(to_unsigned(26, 8)),
			2825 => std_logic_vector(to_unsigned(134, 8)),
			2826 => std_logic_vector(to_unsigned(118, 8)),
			2827 => std_logic_vector(to_unsigned(41, 8)),
			2828 => std_logic_vector(to_unsigned(33, 8)),
			2829 => std_logic_vector(to_unsigned(130, 8)),
			2830 => std_logic_vector(to_unsigned(131, 8)),
			2831 => std_logic_vector(to_unsigned(8, 8)),
			2832 => std_logic_vector(to_unsigned(49, 8)),
			2833 => std_logic_vector(to_unsigned(245, 8)),
			2834 => std_logic_vector(to_unsigned(236, 8)),
			2835 => std_logic_vector(to_unsigned(104, 8)),
			2836 => std_logic_vector(to_unsigned(193, 8)),
			2837 => std_logic_vector(to_unsigned(173, 8)),
			2838 => std_logic_vector(to_unsigned(52, 8)),
			2839 => std_logic_vector(to_unsigned(43, 8)),
			2840 => std_logic_vector(to_unsigned(220, 8)),
			2841 => std_logic_vector(to_unsigned(88, 8)),
			2842 => std_logic_vector(to_unsigned(165, 8)),
			2843 => std_logic_vector(to_unsigned(246, 8)),
			2844 => std_logic_vector(to_unsigned(93, 8)),
			2845 => std_logic_vector(to_unsigned(6, 8)),
			2846 => std_logic_vector(to_unsigned(228, 8)),
			2847 => std_logic_vector(to_unsigned(127, 8)),
			2848 => std_logic_vector(to_unsigned(236, 8)),
			2849 => std_logic_vector(to_unsigned(73, 8)),
			2850 => std_logic_vector(to_unsigned(252, 8)),
			2851 => std_logic_vector(to_unsigned(90, 8)),
			2852 => std_logic_vector(to_unsigned(205, 8)),
			2853 => std_logic_vector(to_unsigned(195, 8)),
			2854 => std_logic_vector(to_unsigned(16, 8)),
			2855 => std_logic_vector(to_unsigned(138, 8)),
			2856 => std_logic_vector(to_unsigned(20, 8)),
			2857 => std_logic_vector(to_unsigned(133, 8)),
			2858 => std_logic_vector(to_unsigned(52, 8)),
			2859 => std_logic_vector(to_unsigned(246, 8)),
			2860 => std_logic_vector(to_unsigned(130, 8)),
			2861 => std_logic_vector(to_unsigned(136, 8)),
			2862 => std_logic_vector(to_unsigned(237, 8)),
			2863 => std_logic_vector(to_unsigned(181, 8)),
			2864 => std_logic_vector(to_unsigned(215, 8)),
			2865 => std_logic_vector(to_unsigned(9, 8)),
			2866 => std_logic_vector(to_unsigned(90, 8)),
			2867 => std_logic_vector(to_unsigned(137, 8)),
			2868 => std_logic_vector(to_unsigned(88, 8)),
			2869 => std_logic_vector(to_unsigned(175, 8)),
			2870 => std_logic_vector(to_unsigned(154, 8)),
			2871 => std_logic_vector(to_unsigned(165, 8)),
			2872 => std_logic_vector(to_unsigned(238, 8)),
			2873 => std_logic_vector(to_unsigned(42, 8)),
			2874 => std_logic_vector(to_unsigned(114, 8)),
			2875 => std_logic_vector(to_unsigned(245, 8)),
			2876 => std_logic_vector(to_unsigned(8, 8)),
			2877 => std_logic_vector(to_unsigned(195, 8)),
			2878 => std_logic_vector(to_unsigned(37, 8)),
			2879 => std_logic_vector(to_unsigned(229, 8)),
			2880 => std_logic_vector(to_unsigned(162, 8)),
			2881 => std_logic_vector(to_unsigned(34, 8)),
			2882 => std_logic_vector(to_unsigned(208, 8)),
			2883 => std_logic_vector(to_unsigned(111, 8)),
			2884 => std_logic_vector(to_unsigned(29, 8)),
			2885 => std_logic_vector(to_unsigned(197, 8)),
			2886 => std_logic_vector(to_unsigned(194, 8)),
			2887 => std_logic_vector(to_unsigned(216, 8)),
			2888 => std_logic_vector(to_unsigned(119, 8)),
			2889 => std_logic_vector(to_unsigned(55, 8)),
			2890 => std_logic_vector(to_unsigned(139, 8)),
			2891 => std_logic_vector(to_unsigned(185, 8)),
			2892 => std_logic_vector(to_unsigned(221, 8)),
			2893 => std_logic_vector(to_unsigned(102, 8)),
			2894 => std_logic_vector(to_unsigned(29, 8)),
			2895 => std_logic_vector(to_unsigned(26, 8)),
			2896 => std_logic_vector(to_unsigned(107, 8)),
			2897 => std_logic_vector(to_unsigned(47, 8)),
			2898 => std_logic_vector(to_unsigned(40, 8)),
			2899 => std_logic_vector(to_unsigned(236, 8)),
			2900 => std_logic_vector(to_unsigned(194, 8)),
			2901 => std_logic_vector(to_unsigned(99, 8)),
			2902 => std_logic_vector(to_unsigned(128, 8)),
			2903 => std_logic_vector(to_unsigned(209, 8)),
			2904 => std_logic_vector(to_unsigned(109, 8)),
			2905 => std_logic_vector(to_unsigned(250, 8)),
			2906 => std_logic_vector(to_unsigned(236, 8)),
			2907 => std_logic_vector(to_unsigned(190, 8)),
			2908 => std_logic_vector(to_unsigned(118, 8)),
			2909 => std_logic_vector(to_unsigned(71, 8)),
			2910 => std_logic_vector(to_unsigned(94, 8)),
			2911 => std_logic_vector(to_unsigned(138, 8)),
			2912 => std_logic_vector(to_unsigned(206, 8)),
			2913 => std_logic_vector(to_unsigned(219, 8)),
			2914 => std_logic_vector(to_unsigned(54, 8)),
			2915 => std_logic_vector(to_unsigned(190, 8)),
			2916 => std_logic_vector(to_unsigned(142, 8)),
			2917 => std_logic_vector(to_unsigned(187, 8)),
			2918 => std_logic_vector(to_unsigned(154, 8)),
			2919 => std_logic_vector(to_unsigned(218, 8)),
			2920 => std_logic_vector(to_unsigned(203, 8)),
			2921 => std_logic_vector(to_unsigned(130, 8)),
			2922 => std_logic_vector(to_unsigned(22, 8)),
			2923 => std_logic_vector(to_unsigned(179, 8)),
			2924 => std_logic_vector(to_unsigned(68, 8)),
			2925 => std_logic_vector(to_unsigned(126, 8)),
			2926 => std_logic_vector(to_unsigned(149, 8)),
			2927 => std_logic_vector(to_unsigned(239, 8)),
			2928 => std_logic_vector(to_unsigned(61, 8)),
			2929 => std_logic_vector(to_unsigned(13, 8)),
			2930 => std_logic_vector(to_unsigned(160, 8)),
			2931 => std_logic_vector(to_unsigned(47, 8)),
			2932 => std_logic_vector(to_unsigned(19, 8)),
			2933 => std_logic_vector(to_unsigned(21, 8)),
			2934 => std_logic_vector(to_unsigned(90, 8)),
			2935 => std_logic_vector(to_unsigned(112, 8)),
			2936 => std_logic_vector(to_unsigned(14, 8)),
			2937 => std_logic_vector(to_unsigned(176, 8)),
			2938 => std_logic_vector(to_unsigned(113, 8)),
			2939 => std_logic_vector(to_unsigned(0, 8)),
			2940 => std_logic_vector(to_unsigned(140, 8)),
			2941 => std_logic_vector(to_unsigned(250, 8)),
			2942 => std_logic_vector(to_unsigned(253, 8)),
			2943 => std_logic_vector(to_unsigned(42, 8)),
			2944 => std_logic_vector(to_unsigned(49, 8)),
			2945 => std_logic_vector(to_unsigned(5, 8)),
			2946 => std_logic_vector(to_unsigned(215, 8)),
			2947 => std_logic_vector(to_unsigned(228, 8)),
			2948 => std_logic_vector(to_unsigned(192, 8)),
			2949 => std_logic_vector(to_unsigned(13, 8)),
			2950 => std_logic_vector(to_unsigned(162, 8)),
			2951 => std_logic_vector(to_unsigned(215, 8)),
			2952 => std_logic_vector(to_unsigned(27, 8)),
			2953 => std_logic_vector(to_unsigned(206, 8)),
			2954 => std_logic_vector(to_unsigned(197, 8)),
			2955 => std_logic_vector(to_unsigned(27, 8)),
			2956 => std_logic_vector(to_unsigned(35, 8)),
			2957 => std_logic_vector(to_unsigned(194, 8)),
			2958 => std_logic_vector(to_unsigned(3, 8)),
			2959 => std_logic_vector(to_unsigned(123, 8)),
			2960 => std_logic_vector(to_unsigned(161, 8)),
			2961 => std_logic_vector(to_unsigned(196, 8)),
			2962 => std_logic_vector(to_unsigned(211, 8)),
			2963 => std_logic_vector(to_unsigned(102, 8)),
			2964 => std_logic_vector(to_unsigned(35, 8)),
			2965 => std_logic_vector(to_unsigned(72, 8)),
			2966 => std_logic_vector(to_unsigned(50, 8)),
			2967 => std_logic_vector(to_unsigned(250, 8)),
			2968 => std_logic_vector(to_unsigned(226, 8)),
			2969 => std_logic_vector(to_unsigned(120, 8)),
			2970 => std_logic_vector(to_unsigned(94, 8)),
			2971 => std_logic_vector(to_unsigned(224, 8)),
			2972 => std_logic_vector(to_unsigned(136, 8)),
			2973 => std_logic_vector(to_unsigned(221, 8)),
			2974 => std_logic_vector(to_unsigned(16, 8)),
			2975 => std_logic_vector(to_unsigned(141, 8)),
			2976 => std_logic_vector(to_unsigned(228, 8)),
			2977 => std_logic_vector(to_unsigned(193, 8)),
			2978 => std_logic_vector(to_unsigned(167, 8)),
			2979 => std_logic_vector(to_unsigned(32, 8)),
			2980 => std_logic_vector(to_unsigned(163, 8)),
			2981 => std_logic_vector(to_unsigned(139, 8)),
			2982 => std_logic_vector(to_unsigned(3, 8)),
			2983 => std_logic_vector(to_unsigned(158, 8)),
			2984 => std_logic_vector(to_unsigned(140, 8)),
			2985 => std_logic_vector(to_unsigned(212, 8)),
			2986 => std_logic_vector(to_unsigned(111, 8)),
			2987 => std_logic_vector(to_unsigned(129, 8)),
			2988 => std_logic_vector(to_unsigned(122, 8)),
			2989 => std_logic_vector(to_unsigned(167, 8)),
			2990 => std_logic_vector(to_unsigned(119, 8)),
			2991 => std_logic_vector(to_unsigned(99, 8)),
			2992 => std_logic_vector(to_unsigned(82, 8)),
			2993 => std_logic_vector(to_unsigned(238, 8)),
			2994 => std_logic_vector(to_unsigned(139, 8)),
			2995 => std_logic_vector(to_unsigned(81, 8)),
			2996 => std_logic_vector(to_unsigned(79, 8)),
			2997 => std_logic_vector(to_unsigned(26, 8)),
			2998 => std_logic_vector(to_unsigned(200, 8)),
			2999 => std_logic_vector(to_unsigned(5, 8)),
			3000 => std_logic_vector(to_unsigned(109, 8)),
			3001 => std_logic_vector(to_unsigned(109, 8)),
			3002 => std_logic_vector(to_unsigned(55, 8)),
			3003 => std_logic_vector(to_unsigned(176, 8)),
			3004 => std_logic_vector(to_unsigned(158, 8)),
			3005 => std_logic_vector(to_unsigned(152, 8)),
			3006 => std_logic_vector(to_unsigned(251, 8)),
			3007 => std_logic_vector(to_unsigned(250, 8)),
			3008 => std_logic_vector(to_unsigned(81, 8)),
			3009 => std_logic_vector(to_unsigned(15, 8)),
			3010 => std_logic_vector(to_unsigned(139, 8)),
			3011 => std_logic_vector(to_unsigned(158, 8)),
			3012 => std_logic_vector(to_unsigned(173, 8)),
			3013 => std_logic_vector(to_unsigned(74, 8)),
			3014 => std_logic_vector(to_unsigned(245, 8)),
			3015 => std_logic_vector(to_unsigned(149, 8)),
			3016 => std_logic_vector(to_unsigned(80, 8)),
			3017 => std_logic_vector(to_unsigned(210, 8)),
			3018 => std_logic_vector(to_unsigned(33, 8)),
			3019 => std_logic_vector(to_unsigned(207, 8)),
			3020 => std_logic_vector(to_unsigned(9, 8)),
			3021 => std_logic_vector(to_unsigned(228, 8)),
			3022 => std_logic_vector(to_unsigned(251, 8)),
			3023 => std_logic_vector(to_unsigned(38, 8)),
			3024 => std_logic_vector(to_unsigned(87, 8)),
			3025 => std_logic_vector(to_unsigned(255, 8)),
			3026 => std_logic_vector(to_unsigned(54, 8)),
			3027 => std_logic_vector(to_unsigned(85, 8)),
			3028 => std_logic_vector(to_unsigned(98, 8)),
			3029 => std_logic_vector(to_unsigned(10, 8)),
			3030 => std_logic_vector(to_unsigned(128, 8)),
			3031 => std_logic_vector(to_unsigned(59, 8)),
			3032 => std_logic_vector(to_unsigned(28, 8)),
			3033 => std_logic_vector(to_unsigned(57, 8)),
			3034 => std_logic_vector(to_unsigned(163, 8)),
			3035 => std_logic_vector(to_unsigned(95, 8)),
			3036 => std_logic_vector(to_unsigned(25, 8)),
			3037 => std_logic_vector(to_unsigned(62, 8)),
			3038 => std_logic_vector(to_unsigned(148, 8)),
			3039 => std_logic_vector(to_unsigned(48, 8)),
			3040 => std_logic_vector(to_unsigned(163, 8)),
			3041 => std_logic_vector(to_unsigned(84, 8)),
			3042 => std_logic_vector(to_unsigned(225, 8)),
			3043 => std_logic_vector(to_unsigned(225, 8)),
			3044 => std_logic_vector(to_unsigned(163, 8)),
			3045 => std_logic_vector(to_unsigned(174, 8)),
			3046 => std_logic_vector(to_unsigned(63, 8)),
			3047 => std_logic_vector(to_unsigned(85, 8)),
			3048 => std_logic_vector(to_unsigned(152, 8)),
			3049 => std_logic_vector(to_unsigned(233, 8)),
			3050 => std_logic_vector(to_unsigned(66, 8)),
			3051 => std_logic_vector(to_unsigned(240, 8)),
			3052 => std_logic_vector(to_unsigned(255, 8)),
			3053 => std_logic_vector(to_unsigned(88, 8)),
			3054 => std_logic_vector(to_unsigned(15, 8)),
			3055 => std_logic_vector(to_unsigned(114, 8)),
			3056 => std_logic_vector(to_unsigned(190, 8)),
			3057 => std_logic_vector(to_unsigned(111, 8)),
			3058 => std_logic_vector(to_unsigned(12, 8)),
			3059 => std_logic_vector(to_unsigned(166, 8)),
			3060 => std_logic_vector(to_unsigned(167, 8)),
			3061 => std_logic_vector(to_unsigned(41, 8)),
			3062 => std_logic_vector(to_unsigned(107, 8)),
			3063 => std_logic_vector(to_unsigned(117, 8)),
			3064 => std_logic_vector(to_unsigned(114, 8)),
			3065 => std_logic_vector(to_unsigned(62, 8)),
			3066 => std_logic_vector(to_unsigned(74, 8)),
			3067 => std_logic_vector(to_unsigned(94, 8)),
			3068 => std_logic_vector(to_unsigned(205, 8)),
			3069 => std_logic_vector(to_unsigned(195, 8)),
			3070 => std_logic_vector(to_unsigned(43, 8)),
			3071 => std_logic_vector(to_unsigned(37, 8)),
			3072 => std_logic_vector(to_unsigned(246, 8)),
			3073 => std_logic_vector(to_unsigned(0, 8)),
			3074 => std_logic_vector(to_unsigned(141, 8)),
			3075 => std_logic_vector(to_unsigned(203, 8)),
			3076 => std_logic_vector(to_unsigned(100, 8)),
			3077 => std_logic_vector(to_unsigned(231, 8)),
			3078 => std_logic_vector(to_unsigned(89, 8)),
			3079 => std_logic_vector(to_unsigned(89, 8)),
			3080 => std_logic_vector(to_unsigned(169, 8)),
			3081 => std_logic_vector(to_unsigned(190, 8)),
			3082 => std_logic_vector(to_unsigned(167, 8)),
			3083 => std_logic_vector(to_unsigned(194, 8)),
			3084 => std_logic_vector(to_unsigned(63, 8)),
			3085 => std_logic_vector(to_unsigned(18, 8)),
			3086 => std_logic_vector(to_unsigned(224, 8)),
			3087 => std_logic_vector(to_unsigned(41, 8)),
			3088 => std_logic_vector(to_unsigned(100, 8)),
			3089 => std_logic_vector(to_unsigned(97, 8)),
			3090 => std_logic_vector(to_unsigned(54, 8)),
			3091 => std_logic_vector(to_unsigned(172, 8)),
			3092 => std_logic_vector(to_unsigned(10, 8)),
			3093 => std_logic_vector(to_unsigned(127, 8)),
			3094 => std_logic_vector(to_unsigned(233, 8)),
			3095 => std_logic_vector(to_unsigned(4, 8)),
			3096 => std_logic_vector(to_unsigned(126, 8)),
			3097 => std_logic_vector(to_unsigned(86, 8)),
			3098 => std_logic_vector(to_unsigned(108, 8)),
			3099 => std_logic_vector(to_unsigned(123, 8)),
			3100 => std_logic_vector(to_unsigned(161, 8)),
			3101 => std_logic_vector(to_unsigned(236, 8)),
			3102 => std_logic_vector(to_unsigned(153, 8)),
			3103 => std_logic_vector(to_unsigned(132, 8)),
			3104 => std_logic_vector(to_unsigned(215, 8)),
			3105 => std_logic_vector(to_unsigned(140, 8)),
			3106 => std_logic_vector(to_unsigned(30, 8)),
			3107 => std_logic_vector(to_unsigned(5, 8)),
			3108 => std_logic_vector(to_unsigned(113, 8)),
			3109 => std_logic_vector(to_unsigned(9, 8)),
			3110 => std_logic_vector(to_unsigned(236, 8)),
			3111 => std_logic_vector(to_unsigned(138, 8)),
			3112 => std_logic_vector(to_unsigned(34, 8)),
			3113 => std_logic_vector(to_unsigned(152, 8)),
			3114 => std_logic_vector(to_unsigned(141, 8)),
			3115 => std_logic_vector(to_unsigned(169, 8)),
			3116 => std_logic_vector(to_unsigned(57, 8)),
			3117 => std_logic_vector(to_unsigned(86, 8)),
			3118 => std_logic_vector(to_unsigned(88, 8)),
			3119 => std_logic_vector(to_unsigned(235, 8)),
			3120 => std_logic_vector(to_unsigned(33, 8)),
			3121 => std_logic_vector(to_unsigned(186, 8)),
			3122 => std_logic_vector(to_unsigned(86, 8)),
			3123 => std_logic_vector(to_unsigned(42, 8)),
			3124 => std_logic_vector(to_unsigned(121, 8)),
			3125 => std_logic_vector(to_unsigned(108, 8)),
			3126 => std_logic_vector(to_unsigned(207, 8)),
			3127 => std_logic_vector(to_unsigned(245, 8)),
			3128 => std_logic_vector(to_unsigned(243, 8)),
			3129 => std_logic_vector(to_unsigned(174, 8)),
			3130 => std_logic_vector(to_unsigned(139, 8)),
			3131 => std_logic_vector(to_unsigned(200, 8)),
			3132 => std_logic_vector(to_unsigned(70, 8)),
			3133 => std_logic_vector(to_unsigned(143, 8)),
			3134 => std_logic_vector(to_unsigned(135, 8)),
			3135 => std_logic_vector(to_unsigned(229, 8)),
			3136 => std_logic_vector(to_unsigned(216, 8)),
			3137 => std_logic_vector(to_unsigned(36, 8)),
			3138 => std_logic_vector(to_unsigned(42, 8)),
			3139 => std_logic_vector(to_unsigned(117, 8)),
			3140 => std_logic_vector(to_unsigned(204, 8)),
			3141 => std_logic_vector(to_unsigned(203, 8)),
			3142 => std_logic_vector(to_unsigned(27, 8)),
			3143 => std_logic_vector(to_unsigned(178, 8)),
			3144 => std_logic_vector(to_unsigned(106, 8)),
			3145 => std_logic_vector(to_unsigned(74, 8)),
			3146 => std_logic_vector(to_unsigned(195, 8)),
			3147 => std_logic_vector(to_unsigned(128, 8)),
			3148 => std_logic_vector(to_unsigned(223, 8)),
			3149 => std_logic_vector(to_unsigned(178, 8)),
			3150 => std_logic_vector(to_unsigned(170, 8)),
			3151 => std_logic_vector(to_unsigned(231, 8)),
			3152 => std_logic_vector(to_unsigned(213, 8)),
			3153 => std_logic_vector(to_unsigned(146, 8)),
			3154 => std_logic_vector(to_unsigned(24, 8)),
			3155 => std_logic_vector(to_unsigned(119, 8)),
			3156 => std_logic_vector(to_unsigned(182, 8)),
			3157 => std_logic_vector(to_unsigned(100, 8)),
			3158 => std_logic_vector(to_unsigned(142, 8)),
			3159 => std_logic_vector(to_unsigned(149, 8)),
			3160 => std_logic_vector(to_unsigned(125, 8)),
			3161 => std_logic_vector(to_unsigned(246, 8)),
			3162 => std_logic_vector(to_unsigned(152, 8)),
			3163 => std_logic_vector(to_unsigned(11, 8)),
			3164 => std_logic_vector(to_unsigned(34, 8)),
			3165 => std_logic_vector(to_unsigned(178, 8)),
			3166 => std_logic_vector(to_unsigned(25, 8)),
			3167 => std_logic_vector(to_unsigned(185, 8)),
			3168 => std_logic_vector(to_unsigned(54, 8)),
			3169 => std_logic_vector(to_unsigned(248, 8)),
			3170 => std_logic_vector(to_unsigned(92, 8)),
			3171 => std_logic_vector(to_unsigned(218, 8)),
			3172 => std_logic_vector(to_unsigned(132, 8)),
			3173 => std_logic_vector(to_unsigned(20, 8)),
			3174 => std_logic_vector(to_unsigned(223, 8)),
			3175 => std_logic_vector(to_unsigned(214, 8)),
			3176 => std_logic_vector(to_unsigned(38, 8)),
			3177 => std_logic_vector(to_unsigned(130, 8)),
			3178 => std_logic_vector(to_unsigned(114, 8)),
			3179 => std_logic_vector(to_unsigned(218, 8)),
			3180 => std_logic_vector(to_unsigned(206, 8)),
			3181 => std_logic_vector(to_unsigned(229, 8)),
			3182 => std_logic_vector(to_unsigned(204, 8)),
			3183 => std_logic_vector(to_unsigned(141, 8)),
			3184 => std_logic_vector(to_unsigned(160, 8)),
			3185 => std_logic_vector(to_unsigned(104, 8)),
			3186 => std_logic_vector(to_unsigned(187, 8)),
			3187 => std_logic_vector(to_unsigned(112, 8)),
			3188 => std_logic_vector(to_unsigned(201, 8)),
			3189 => std_logic_vector(to_unsigned(26, 8)),
			3190 => std_logic_vector(to_unsigned(165, 8)),
			3191 => std_logic_vector(to_unsigned(139, 8)),
			3192 => std_logic_vector(to_unsigned(103, 8)),
			3193 => std_logic_vector(to_unsigned(127, 8)),
			3194 => std_logic_vector(to_unsigned(99, 8)),
			3195 => std_logic_vector(to_unsigned(183, 8)),
			3196 => std_logic_vector(to_unsigned(3, 8)),
			3197 => std_logic_vector(to_unsigned(125, 8)),
			3198 => std_logic_vector(to_unsigned(192, 8)),
			3199 => std_logic_vector(to_unsigned(229, 8)),
			3200 => std_logic_vector(to_unsigned(136, 8)),
			3201 => std_logic_vector(to_unsigned(63, 8)),
			3202 => std_logic_vector(to_unsigned(18, 8)),
			3203 => std_logic_vector(to_unsigned(170, 8)),
			3204 => std_logic_vector(to_unsigned(117, 8)),
			3205 => std_logic_vector(to_unsigned(130, 8)),
			3206 => std_logic_vector(to_unsigned(223, 8)),
			3207 => std_logic_vector(to_unsigned(104, 8)),
			3208 => std_logic_vector(to_unsigned(202, 8)),
			3209 => std_logic_vector(to_unsigned(16, 8)),
			3210 => std_logic_vector(to_unsigned(101, 8)),
			3211 => std_logic_vector(to_unsigned(52, 8)),
			3212 => std_logic_vector(to_unsigned(234, 8)),
			3213 => std_logic_vector(to_unsigned(14, 8)),
			3214 => std_logic_vector(to_unsigned(9, 8)),
			3215 => std_logic_vector(to_unsigned(221, 8)),
			3216 => std_logic_vector(to_unsigned(6, 8)),
			3217 => std_logic_vector(to_unsigned(166, 8)),
			3218 => std_logic_vector(to_unsigned(160, 8)),
			3219 => std_logic_vector(to_unsigned(200, 8)),
			3220 => std_logic_vector(to_unsigned(217, 8)),
			3221 => std_logic_vector(to_unsigned(216, 8)),
			3222 => std_logic_vector(to_unsigned(172, 8)),
			3223 => std_logic_vector(to_unsigned(243, 8)),
			3224 => std_logic_vector(to_unsigned(10, 8)),
			3225 => std_logic_vector(to_unsigned(184, 8)),
			3226 => std_logic_vector(to_unsigned(220, 8)),
			3227 => std_logic_vector(to_unsigned(69, 8)),
			3228 => std_logic_vector(to_unsigned(116, 8)),
			3229 => std_logic_vector(to_unsigned(147, 8)),
			3230 => std_logic_vector(to_unsigned(212, 8)),
			3231 => std_logic_vector(to_unsigned(185, 8)),
			3232 => std_logic_vector(to_unsigned(3, 8)),
			3233 => std_logic_vector(to_unsigned(155, 8)),
			3234 => std_logic_vector(to_unsigned(175, 8)),
			3235 => std_logic_vector(to_unsigned(46, 8)),
			3236 => std_logic_vector(to_unsigned(221, 8)),
			3237 => std_logic_vector(to_unsigned(240, 8)),
			3238 => std_logic_vector(to_unsigned(250, 8)),
			3239 => std_logic_vector(to_unsigned(5, 8)),
			3240 => std_logic_vector(to_unsigned(85, 8)),
			3241 => std_logic_vector(to_unsigned(95, 8)),
			3242 => std_logic_vector(to_unsigned(92, 8)),
			3243 => std_logic_vector(to_unsigned(42, 8)),
			3244 => std_logic_vector(to_unsigned(84, 8)),
			3245 => std_logic_vector(to_unsigned(138, 8)),
			3246 => std_logic_vector(to_unsigned(138, 8)),
			3247 => std_logic_vector(to_unsigned(172, 8)),
			3248 => std_logic_vector(to_unsigned(135, 8)),
			3249 => std_logic_vector(to_unsigned(18, 8)),
			3250 => std_logic_vector(to_unsigned(36, 8)),
			3251 => std_logic_vector(to_unsigned(248, 8)),
			3252 => std_logic_vector(to_unsigned(254, 8)),
			3253 => std_logic_vector(to_unsigned(119, 8)),
			3254 => std_logic_vector(to_unsigned(113, 8)),
			3255 => std_logic_vector(to_unsigned(118, 8)),
			3256 => std_logic_vector(to_unsigned(1, 8)),
			3257 => std_logic_vector(to_unsigned(25, 8)),
			3258 => std_logic_vector(to_unsigned(255, 8)),
			3259 => std_logic_vector(to_unsigned(41, 8)),
			3260 => std_logic_vector(to_unsigned(70, 8)),
			3261 => std_logic_vector(to_unsigned(203, 8)),
			3262 => std_logic_vector(to_unsigned(253, 8)),
			3263 => std_logic_vector(to_unsigned(84, 8)),
			3264 => std_logic_vector(to_unsigned(88, 8)),
			3265 => std_logic_vector(to_unsigned(49, 8)),
			3266 => std_logic_vector(to_unsigned(59, 8)),
			3267 => std_logic_vector(to_unsigned(31, 8)),
			3268 => std_logic_vector(to_unsigned(23, 8)),
			3269 => std_logic_vector(to_unsigned(134, 8)),
			3270 => std_logic_vector(to_unsigned(89, 8)),
			3271 => std_logic_vector(to_unsigned(72, 8)),
			3272 => std_logic_vector(to_unsigned(50, 8)),
			3273 => std_logic_vector(to_unsigned(5, 8)),
			3274 => std_logic_vector(to_unsigned(118, 8)),
			3275 => std_logic_vector(to_unsigned(174, 8)),
			3276 => std_logic_vector(to_unsigned(56, 8)),
			3277 => std_logic_vector(to_unsigned(68, 8)),
			3278 => std_logic_vector(to_unsigned(156, 8)),
			3279 => std_logic_vector(to_unsigned(179, 8)),
			3280 => std_logic_vector(to_unsigned(95, 8)),
			3281 => std_logic_vector(to_unsigned(133, 8)),
			3282 => std_logic_vector(to_unsigned(139, 8)),
			3283 => std_logic_vector(to_unsigned(215, 8)),
			3284 => std_logic_vector(to_unsigned(0, 8)),
			3285 => std_logic_vector(to_unsigned(156, 8)),
			3286 => std_logic_vector(to_unsigned(58, 8)),
			3287 => std_logic_vector(to_unsigned(130, 8)),
			3288 => std_logic_vector(to_unsigned(19, 8)),
			3289 => std_logic_vector(to_unsigned(204, 8)),
			3290 => std_logic_vector(to_unsigned(227, 8)),
			3291 => std_logic_vector(to_unsigned(218, 8)),
			3292 => std_logic_vector(to_unsigned(106, 8)),
			3293 => std_logic_vector(to_unsigned(34, 8)),
			3294 => std_logic_vector(to_unsigned(1, 8)),
			3295 => std_logic_vector(to_unsigned(150, 8)),
			3296 => std_logic_vector(to_unsigned(249, 8)),
			3297 => std_logic_vector(to_unsigned(101, 8)),
			3298 => std_logic_vector(to_unsigned(224, 8)),
			3299 => std_logic_vector(to_unsigned(113, 8)),
			3300 => std_logic_vector(to_unsigned(159, 8)),
			3301 => std_logic_vector(to_unsigned(201, 8)),
			3302 => std_logic_vector(to_unsigned(28, 8)),
			3303 => std_logic_vector(to_unsigned(116, 8)),
			3304 => std_logic_vector(to_unsigned(33, 8)),
			3305 => std_logic_vector(to_unsigned(193, 8)),
			3306 => std_logic_vector(to_unsigned(153, 8)),
			3307 => std_logic_vector(to_unsigned(222, 8)),
			3308 => std_logic_vector(to_unsigned(221, 8)),
			3309 => std_logic_vector(to_unsigned(172, 8)),
			3310 => std_logic_vector(to_unsigned(126, 8)),
			3311 => std_logic_vector(to_unsigned(192, 8)),
			3312 => std_logic_vector(to_unsigned(116, 8)),
			3313 => std_logic_vector(to_unsigned(48, 8)),
			3314 => std_logic_vector(to_unsigned(136, 8)),
			3315 => std_logic_vector(to_unsigned(171, 8)),
			3316 => std_logic_vector(to_unsigned(84, 8)),
			3317 => std_logic_vector(to_unsigned(71, 8)),
			3318 => std_logic_vector(to_unsigned(105, 8)),
			3319 => std_logic_vector(to_unsigned(46, 8)),
			3320 => std_logic_vector(to_unsigned(127, 8)),
			3321 => std_logic_vector(to_unsigned(242, 8)),
			3322 => std_logic_vector(to_unsigned(54, 8)),
			3323 => std_logic_vector(to_unsigned(81, 8)),
			3324 => std_logic_vector(to_unsigned(201, 8)),
			3325 => std_logic_vector(to_unsigned(196, 8)),
			3326 => std_logic_vector(to_unsigned(170, 8)),
			3327 => std_logic_vector(to_unsigned(120, 8)),
			3328 => std_logic_vector(to_unsigned(87, 8)),
			3329 => std_logic_vector(to_unsigned(64, 8)),
			3330 => std_logic_vector(to_unsigned(197, 8)),
			3331 => std_logic_vector(to_unsigned(56, 8)),
			3332 => std_logic_vector(to_unsigned(248, 8)),
			3333 => std_logic_vector(to_unsigned(66, 8)),
			3334 => std_logic_vector(to_unsigned(49, 8)),
			3335 => std_logic_vector(to_unsigned(237, 8)),
			3336 => std_logic_vector(to_unsigned(74, 8)),
			3337 => std_logic_vector(to_unsigned(79, 8)),
			3338 => std_logic_vector(to_unsigned(141, 8)),
			3339 => std_logic_vector(to_unsigned(27, 8)),
			3340 => std_logic_vector(to_unsigned(180, 8)),
			3341 => std_logic_vector(to_unsigned(120, 8)),
			3342 => std_logic_vector(to_unsigned(157, 8)),
			3343 => std_logic_vector(to_unsigned(122, 8)),
			3344 => std_logic_vector(to_unsigned(18, 8)),
			3345 => std_logic_vector(to_unsigned(85, 8)),
			3346 => std_logic_vector(to_unsigned(224, 8)),
			3347 => std_logic_vector(to_unsigned(81, 8)),
			3348 => std_logic_vector(to_unsigned(185, 8)),
			3349 => std_logic_vector(to_unsigned(175, 8)),
			3350 => std_logic_vector(to_unsigned(205, 8)),
			3351 => std_logic_vector(to_unsigned(18, 8)),
			3352 => std_logic_vector(to_unsigned(9, 8)),
			3353 => std_logic_vector(to_unsigned(89, 8)),
			3354 => std_logic_vector(to_unsigned(201, 8)),
			3355 => std_logic_vector(to_unsigned(91, 8)),
			3356 => std_logic_vector(to_unsigned(162, 8)),
			3357 => std_logic_vector(to_unsigned(14, 8)),
			3358 => std_logic_vector(to_unsigned(76, 8)),
			3359 => std_logic_vector(to_unsigned(74, 8)),
			3360 => std_logic_vector(to_unsigned(94, 8)),
			3361 => std_logic_vector(to_unsigned(71, 8)),
			3362 => std_logic_vector(to_unsigned(175, 8)),
			3363 => std_logic_vector(to_unsigned(192, 8)),
			3364 => std_logic_vector(to_unsigned(137, 8)),
			3365 => std_logic_vector(to_unsigned(134, 8)),
			3366 => std_logic_vector(to_unsigned(180, 8)),
			3367 => std_logic_vector(to_unsigned(213, 8)),
			3368 => std_logic_vector(to_unsigned(174, 8)),
			3369 => std_logic_vector(to_unsigned(205, 8)),
			3370 => std_logic_vector(to_unsigned(163, 8)),
			3371 => std_logic_vector(to_unsigned(111, 8)),
			3372 => std_logic_vector(to_unsigned(129, 8)),
			3373 => std_logic_vector(to_unsigned(1, 8)),
			3374 => std_logic_vector(to_unsigned(40, 8)),
			3375 => std_logic_vector(to_unsigned(255, 8)),
			3376 => std_logic_vector(to_unsigned(162, 8)),
			3377 => std_logic_vector(to_unsigned(62, 8)),
			3378 => std_logic_vector(to_unsigned(225, 8)),
			3379 => std_logic_vector(to_unsigned(140, 8)),
			3380 => std_logic_vector(to_unsigned(100, 8)),
			3381 => std_logic_vector(to_unsigned(99, 8)),
			3382 => std_logic_vector(to_unsigned(106, 8)),
			3383 => std_logic_vector(to_unsigned(81, 8)),
			3384 => std_logic_vector(to_unsigned(127, 8)),
			3385 => std_logic_vector(to_unsigned(218, 8)),
			3386 => std_logic_vector(to_unsigned(69, 8)),
			3387 => std_logic_vector(to_unsigned(206, 8)),
			3388 => std_logic_vector(to_unsigned(230, 8)),
			3389 => std_logic_vector(to_unsigned(162, 8)),
			3390 => std_logic_vector(to_unsigned(220, 8)),
			3391 => std_logic_vector(to_unsigned(18, 8)),
			3392 => std_logic_vector(to_unsigned(93, 8)),
			3393 => std_logic_vector(to_unsigned(149, 8)),
			3394 => std_logic_vector(to_unsigned(121, 8)),
			3395 => std_logic_vector(to_unsigned(56, 8)),
			3396 => std_logic_vector(to_unsigned(175, 8)),
			3397 => std_logic_vector(to_unsigned(106, 8)),
			3398 => std_logic_vector(to_unsigned(85, 8)),
			3399 => std_logic_vector(to_unsigned(187, 8)),
			3400 => std_logic_vector(to_unsigned(105, 8)),
			3401 => std_logic_vector(to_unsigned(130, 8)),
			3402 => std_logic_vector(to_unsigned(193, 8)),
			3403 => std_logic_vector(to_unsigned(200, 8)),
			3404 => std_logic_vector(to_unsigned(173, 8)),
			3405 => std_logic_vector(to_unsigned(79, 8)),
			3406 => std_logic_vector(to_unsigned(152, 8)),
			3407 => std_logic_vector(to_unsigned(87, 8)),
			3408 => std_logic_vector(to_unsigned(242, 8)),
			3409 => std_logic_vector(to_unsigned(220, 8)),
			3410 => std_logic_vector(to_unsigned(136, 8)),
			3411 => std_logic_vector(to_unsigned(179, 8)),
			3412 => std_logic_vector(to_unsigned(34, 8)),
			3413 => std_logic_vector(to_unsigned(119, 8)),
			3414 => std_logic_vector(to_unsigned(30, 8)),
			3415 => std_logic_vector(to_unsigned(172, 8)),
			3416 => std_logic_vector(to_unsigned(103, 8)),
			3417 => std_logic_vector(to_unsigned(181, 8)),
			3418 => std_logic_vector(to_unsigned(4, 8)),
			3419 => std_logic_vector(to_unsigned(23, 8)),
			3420 => std_logic_vector(to_unsigned(175, 8)),
			3421 => std_logic_vector(to_unsigned(91, 8)),
			3422 => std_logic_vector(to_unsigned(150, 8)),
			3423 => std_logic_vector(to_unsigned(140, 8)),
			3424 => std_logic_vector(to_unsigned(126, 8)),
			3425 => std_logic_vector(to_unsigned(206, 8)),
			3426 => std_logic_vector(to_unsigned(41, 8)),
			3427 => std_logic_vector(to_unsigned(180, 8)),
			3428 => std_logic_vector(to_unsigned(19, 8)),
			3429 => std_logic_vector(to_unsigned(63, 8)),
			3430 => std_logic_vector(to_unsigned(22, 8)),
			3431 => std_logic_vector(to_unsigned(138, 8)),
			3432 => std_logic_vector(to_unsigned(2, 8)),
			3433 => std_logic_vector(to_unsigned(176, 8)),
			3434 => std_logic_vector(to_unsigned(209, 8)),
			3435 => std_logic_vector(to_unsigned(52, 8)),
			3436 => std_logic_vector(to_unsigned(252, 8)),
			3437 => std_logic_vector(to_unsigned(38, 8)),
			3438 => std_logic_vector(to_unsigned(207, 8)),
			3439 => std_logic_vector(to_unsigned(139, 8)),
			3440 => std_logic_vector(to_unsigned(134, 8)),
			3441 => std_logic_vector(to_unsigned(179, 8)),
			3442 => std_logic_vector(to_unsigned(195, 8)),
			3443 => std_logic_vector(to_unsigned(62, 8)),
			3444 => std_logic_vector(to_unsigned(223, 8)),
			3445 => std_logic_vector(to_unsigned(250, 8)),
			3446 => std_logic_vector(to_unsigned(120, 8)),
			3447 => std_logic_vector(to_unsigned(161, 8)),
			3448 => std_logic_vector(to_unsigned(225, 8)),
			3449 => std_logic_vector(to_unsigned(36, 8)),
			3450 => std_logic_vector(to_unsigned(75, 8)),
			3451 => std_logic_vector(to_unsigned(249, 8)),
			3452 => std_logic_vector(to_unsigned(15, 8)),
			3453 => std_logic_vector(to_unsigned(10, 8)),
			3454 => std_logic_vector(to_unsigned(15, 8)),
			3455 => std_logic_vector(to_unsigned(108, 8)),
			3456 => std_logic_vector(to_unsigned(88, 8)),
			3457 => std_logic_vector(to_unsigned(77, 8)),
			3458 => std_logic_vector(to_unsigned(134, 8)),
			3459 => std_logic_vector(to_unsigned(202, 8)),
			3460 => std_logic_vector(to_unsigned(197, 8)),
			3461 => std_logic_vector(to_unsigned(17, 8)),
			3462 => std_logic_vector(to_unsigned(192, 8)),
			3463 => std_logic_vector(to_unsigned(163, 8)),
			3464 => std_logic_vector(to_unsigned(88, 8)),
			3465 => std_logic_vector(to_unsigned(241, 8)),
			3466 => std_logic_vector(to_unsigned(163, 8)),
			3467 => std_logic_vector(to_unsigned(5, 8)),
			3468 => std_logic_vector(to_unsigned(154, 8)),
			3469 => std_logic_vector(to_unsigned(38, 8)),
			3470 => std_logic_vector(to_unsigned(165, 8)),
			3471 => std_logic_vector(to_unsigned(179, 8)),
			3472 => std_logic_vector(to_unsigned(93, 8)),
			3473 => std_logic_vector(to_unsigned(167, 8)),
			3474 => std_logic_vector(to_unsigned(155, 8)),
			3475 => std_logic_vector(to_unsigned(102, 8)),
			3476 => std_logic_vector(to_unsigned(100, 8)),
			3477 => std_logic_vector(to_unsigned(92, 8)),
			3478 => std_logic_vector(to_unsigned(118, 8)),
			3479 => std_logic_vector(to_unsigned(161, 8)),
			3480 => std_logic_vector(to_unsigned(8, 8)),
			3481 => std_logic_vector(to_unsigned(26, 8)),
			3482 => std_logic_vector(to_unsigned(108, 8)),
			3483 => std_logic_vector(to_unsigned(96, 8)),
			3484 => std_logic_vector(to_unsigned(117, 8)),
			3485 => std_logic_vector(to_unsigned(25, 8)),
			3486 => std_logic_vector(to_unsigned(16, 8)),
			3487 => std_logic_vector(to_unsigned(170, 8)),
			3488 => std_logic_vector(to_unsigned(217, 8)),
			3489 => std_logic_vector(to_unsigned(14, 8)),
			3490 => std_logic_vector(to_unsigned(199, 8)),
			3491 => std_logic_vector(to_unsigned(44, 8)),
			3492 => std_logic_vector(to_unsigned(31, 8)),
			3493 => std_logic_vector(to_unsigned(136, 8)),
			3494 => std_logic_vector(to_unsigned(75, 8)),
			3495 => std_logic_vector(to_unsigned(253, 8)),
			3496 => std_logic_vector(to_unsigned(82, 8)),
			3497 => std_logic_vector(to_unsigned(209, 8)),
			3498 => std_logic_vector(to_unsigned(17, 8)),
			3499 => std_logic_vector(to_unsigned(37, 8)),
			3500 => std_logic_vector(to_unsigned(53, 8)),
			3501 => std_logic_vector(to_unsigned(207, 8)),
			3502 => std_logic_vector(to_unsigned(179, 8)),
			3503 => std_logic_vector(to_unsigned(73, 8)),
			3504 => std_logic_vector(to_unsigned(123, 8)),
			3505 => std_logic_vector(to_unsigned(137, 8)),
			3506 => std_logic_vector(to_unsigned(189, 8)),
			3507 => std_logic_vector(to_unsigned(230, 8)),
			3508 => std_logic_vector(to_unsigned(165, 8)),
			3509 => std_logic_vector(to_unsigned(199, 8)),
			3510 => std_logic_vector(to_unsigned(150, 8)),
			3511 => std_logic_vector(to_unsigned(105, 8)),
			3512 => std_logic_vector(to_unsigned(208, 8)),
			3513 => std_logic_vector(to_unsigned(91, 8)),
			3514 => std_logic_vector(to_unsigned(68, 8)),
			3515 => std_logic_vector(to_unsigned(250, 8)),
			3516 => std_logic_vector(to_unsigned(77, 8)),
			3517 => std_logic_vector(to_unsigned(118, 8)),
			3518 => std_logic_vector(to_unsigned(8, 8)),
			3519 => std_logic_vector(to_unsigned(229, 8)),
			3520 => std_logic_vector(to_unsigned(221, 8)),
			3521 => std_logic_vector(to_unsigned(81, 8)),
			3522 => std_logic_vector(to_unsigned(229, 8)),
			3523 => std_logic_vector(to_unsigned(145, 8)),
			3524 => std_logic_vector(to_unsigned(70, 8)),
			3525 => std_logic_vector(to_unsigned(208, 8)),
			3526 => std_logic_vector(to_unsigned(139, 8)),
			3527 => std_logic_vector(to_unsigned(96, 8)),
			3528 => std_logic_vector(to_unsigned(181, 8)),
			3529 => std_logic_vector(to_unsigned(169, 8)),
			3530 => std_logic_vector(to_unsigned(211, 8)),
			3531 => std_logic_vector(to_unsigned(115, 8)),
			3532 => std_logic_vector(to_unsigned(80, 8)),
			3533 => std_logic_vector(to_unsigned(51, 8)),
			3534 => std_logic_vector(to_unsigned(109, 8)),
			3535 => std_logic_vector(to_unsigned(188, 8)),
			3536 => std_logic_vector(to_unsigned(238, 8)),
			3537 => std_logic_vector(to_unsigned(88, 8)),
			3538 => std_logic_vector(to_unsigned(50, 8)),
			3539 => std_logic_vector(to_unsigned(185, 8)),
			3540 => std_logic_vector(to_unsigned(62, 8)),
			3541 => std_logic_vector(to_unsigned(179, 8)),
			3542 => std_logic_vector(to_unsigned(236, 8)),
			3543 => std_logic_vector(to_unsigned(26, 8)),
			3544 => std_logic_vector(to_unsigned(32, 8)),
			3545 => std_logic_vector(to_unsigned(201, 8)),
			3546 => std_logic_vector(to_unsigned(209, 8)),
			3547 => std_logic_vector(to_unsigned(188, 8)),
			3548 => std_logic_vector(to_unsigned(234, 8)),
			3549 => std_logic_vector(to_unsigned(149, 8)),
			3550 => std_logic_vector(to_unsigned(245, 8)),
			3551 => std_logic_vector(to_unsigned(172, 8)),
			3552 => std_logic_vector(to_unsigned(53, 8)),
			3553 => std_logic_vector(to_unsigned(99, 8)),
			3554 => std_logic_vector(to_unsigned(150, 8)),
			3555 => std_logic_vector(to_unsigned(102, 8)),
			3556 => std_logic_vector(to_unsigned(20, 8)),
			3557 => std_logic_vector(to_unsigned(188, 8)),
			3558 => std_logic_vector(to_unsigned(254, 8)),
			3559 => std_logic_vector(to_unsigned(198, 8)),
			3560 => std_logic_vector(to_unsigned(149, 8)),
			3561 => std_logic_vector(to_unsigned(95, 8)),
			3562 => std_logic_vector(to_unsigned(253, 8)),
			3563 => std_logic_vector(to_unsigned(56, 8)),
			3564 => std_logic_vector(to_unsigned(132, 8)),
			3565 => std_logic_vector(to_unsigned(234, 8)),
			3566 => std_logic_vector(to_unsigned(237, 8)),
			3567 => std_logic_vector(to_unsigned(141, 8)),
			3568 => std_logic_vector(to_unsigned(207, 8)),
			3569 => std_logic_vector(to_unsigned(51, 8)),
			3570 => std_logic_vector(to_unsigned(150, 8)),
			3571 => std_logic_vector(to_unsigned(63, 8)),
			3572 => std_logic_vector(to_unsigned(249, 8)),
			3573 => std_logic_vector(to_unsigned(158, 8)),
			3574 => std_logic_vector(to_unsigned(17, 8)),
			3575 => std_logic_vector(to_unsigned(206, 8)),
			3576 => std_logic_vector(to_unsigned(16, 8)),
			3577 => std_logic_vector(to_unsigned(207, 8)),
			3578 => std_logic_vector(to_unsigned(144, 8)),
			3579 => std_logic_vector(to_unsigned(22, 8)),
			3580 => std_logic_vector(to_unsigned(169, 8)),
			3581 => std_logic_vector(to_unsigned(232, 8)),
			3582 => std_logic_vector(to_unsigned(251, 8)),
			3583 => std_logic_vector(to_unsigned(165, 8)),
			3584 => std_logic_vector(to_unsigned(114, 8)),
			3585 => std_logic_vector(to_unsigned(213, 8)),
			3586 => std_logic_vector(to_unsigned(125, 8)),
			3587 => std_logic_vector(to_unsigned(179, 8)),
			3588 => std_logic_vector(to_unsigned(240, 8)),
			3589 => std_logic_vector(to_unsigned(185, 8)),
			3590 => std_logic_vector(to_unsigned(215, 8)),
			3591 => std_logic_vector(to_unsigned(98, 8)),
			3592 => std_logic_vector(to_unsigned(189, 8)),
			3593 => std_logic_vector(to_unsigned(169, 8)),
			3594 => std_logic_vector(to_unsigned(111, 8)),
			3595 => std_logic_vector(to_unsigned(173, 8)),
			3596 => std_logic_vector(to_unsigned(213, 8)),
			3597 => std_logic_vector(to_unsigned(100, 8)),
			3598 => std_logic_vector(to_unsigned(10, 8)),
			3599 => std_logic_vector(to_unsigned(1, 8)),
			3600 => std_logic_vector(to_unsigned(217, 8)),
			3601 => std_logic_vector(to_unsigned(203, 8)),
			3602 => std_logic_vector(to_unsigned(169, 8)),
			3603 => std_logic_vector(to_unsigned(94, 8)),
			3604 => std_logic_vector(to_unsigned(124, 8)),
			3605 => std_logic_vector(to_unsigned(90, 8)),
			3606 => std_logic_vector(to_unsigned(63, 8)),
			3607 => std_logic_vector(to_unsigned(101, 8)),
			3608 => std_logic_vector(to_unsigned(168, 8)),
			3609 => std_logic_vector(to_unsigned(202, 8)),
			3610 => std_logic_vector(to_unsigned(118, 8)),
			3611 => std_logic_vector(to_unsigned(215, 8)),
			3612 => std_logic_vector(to_unsigned(225, 8)),
			3613 => std_logic_vector(to_unsigned(80, 8)),
			3614 => std_logic_vector(to_unsigned(156, 8)),
			3615 => std_logic_vector(to_unsigned(115, 8)),
			3616 => std_logic_vector(to_unsigned(161, 8)),
			3617 => std_logic_vector(to_unsigned(134, 8)),
			3618 => std_logic_vector(to_unsigned(119, 8)),
			3619 => std_logic_vector(to_unsigned(143, 8)),
			3620 => std_logic_vector(to_unsigned(234, 8)),
			3621 => std_logic_vector(to_unsigned(194, 8)),
			3622 => std_logic_vector(to_unsigned(55, 8)),
			3623 => std_logic_vector(to_unsigned(216, 8)),
			3624 => std_logic_vector(to_unsigned(30, 8)),
			3625 => std_logic_vector(to_unsigned(239, 8)),
			3626 => std_logic_vector(to_unsigned(252, 8)),
			3627 => std_logic_vector(to_unsigned(192, 8)),
			3628 => std_logic_vector(to_unsigned(209, 8)),
			3629 => std_logic_vector(to_unsigned(156, 8)),
			3630 => std_logic_vector(to_unsigned(76, 8)),
			3631 => std_logic_vector(to_unsigned(75, 8)),
			3632 => std_logic_vector(to_unsigned(49, 8)),
			3633 => std_logic_vector(to_unsigned(240, 8)),
			3634 => std_logic_vector(to_unsigned(128, 8)),
			3635 => std_logic_vector(to_unsigned(28, 8)),
			3636 => std_logic_vector(to_unsigned(42, 8)),
			3637 => std_logic_vector(to_unsigned(86, 8)),
			3638 => std_logic_vector(to_unsigned(7, 8)),
			3639 => std_logic_vector(to_unsigned(208, 8)),
			3640 => std_logic_vector(to_unsigned(228, 8)),
			3641 => std_logic_vector(to_unsigned(157, 8)),
			3642 => std_logic_vector(to_unsigned(186, 8)),
			3643 => std_logic_vector(to_unsigned(249, 8)),
			3644 => std_logic_vector(to_unsigned(31, 8)),
			3645 => std_logic_vector(to_unsigned(224, 8)),
			3646 => std_logic_vector(to_unsigned(34, 8)),
			3647 => std_logic_vector(to_unsigned(239, 8)),
			3648 => std_logic_vector(to_unsigned(157, 8)),
			3649 => std_logic_vector(to_unsigned(8, 8)),
			3650 => std_logic_vector(to_unsigned(216, 8)),
			3651 => std_logic_vector(to_unsigned(254, 8)),
			3652 => std_logic_vector(to_unsigned(247, 8)),
			3653 => std_logic_vector(to_unsigned(176, 8)),
			3654 => std_logic_vector(to_unsigned(42, 8)),
			3655 => std_logic_vector(to_unsigned(62, 8)),
			3656 => std_logic_vector(to_unsigned(167, 8)),
			3657 => std_logic_vector(to_unsigned(159, 8)),
			3658 => std_logic_vector(to_unsigned(250, 8)),
			3659 => std_logic_vector(to_unsigned(132, 8)),
			3660 => std_logic_vector(to_unsigned(114, 8)),
			3661 => std_logic_vector(to_unsigned(122, 8)),
			3662 => std_logic_vector(to_unsigned(149, 8)),
			3663 => std_logic_vector(to_unsigned(103, 8)),
			3664 => std_logic_vector(to_unsigned(119, 8)),
			3665 => std_logic_vector(to_unsigned(149, 8)),
			3666 => std_logic_vector(to_unsigned(213, 8)),
			3667 => std_logic_vector(to_unsigned(166, 8)),
			3668 => std_logic_vector(to_unsigned(174, 8)),
			3669 => std_logic_vector(to_unsigned(92, 8)),
			3670 => std_logic_vector(to_unsigned(193, 8)),
			3671 => std_logic_vector(to_unsigned(87, 8)),
			3672 => std_logic_vector(to_unsigned(208, 8)),
			3673 => std_logic_vector(to_unsigned(14, 8)),
			3674 => std_logic_vector(to_unsigned(64, 8)),
			3675 => std_logic_vector(to_unsigned(96, 8)),
			3676 => std_logic_vector(to_unsigned(133, 8)),
			3677 => std_logic_vector(to_unsigned(179, 8)),
			3678 => std_logic_vector(to_unsigned(198, 8)),
			3679 => std_logic_vector(to_unsigned(109, 8)),
			3680 => std_logic_vector(to_unsigned(2, 8)),
			3681 => std_logic_vector(to_unsigned(61, 8)),
			3682 => std_logic_vector(to_unsigned(19, 8)),
			3683 => std_logic_vector(to_unsigned(192, 8)),
			3684 => std_logic_vector(to_unsigned(135, 8)),
			3685 => std_logic_vector(to_unsigned(145, 8)),
			3686 => std_logic_vector(to_unsigned(240, 8)),
			3687 => std_logic_vector(to_unsigned(24, 8)),
			3688 => std_logic_vector(to_unsigned(80, 8)),
			3689 => std_logic_vector(to_unsigned(22, 8)),
			3690 => std_logic_vector(to_unsigned(78, 8)),
			3691 => std_logic_vector(to_unsigned(126, 8)),
			3692 => std_logic_vector(to_unsigned(169, 8)),
			3693 => std_logic_vector(to_unsigned(105, 8)),
			3694 => std_logic_vector(to_unsigned(112, 8)),
			3695 => std_logic_vector(to_unsigned(193, 8)),
			3696 => std_logic_vector(to_unsigned(99, 8)),
			3697 => std_logic_vector(to_unsigned(40, 8)),
			3698 => std_logic_vector(to_unsigned(51, 8)),
			3699 => std_logic_vector(to_unsigned(113, 8)),
			3700 => std_logic_vector(to_unsigned(12, 8)),
			3701 => std_logic_vector(to_unsigned(229, 8)),
			3702 => std_logic_vector(to_unsigned(231, 8)),
			3703 => std_logic_vector(to_unsigned(160, 8)),
			3704 => std_logic_vector(to_unsigned(131, 8)),
			3705 => std_logic_vector(to_unsigned(50, 8)),
			3706 => std_logic_vector(to_unsigned(181, 8)),
			3707 => std_logic_vector(to_unsigned(250, 8)),
			3708 => std_logic_vector(to_unsigned(85, 8)),
			3709 => std_logic_vector(to_unsigned(160, 8)),
			3710 => std_logic_vector(to_unsigned(75, 8)),
			3711 => std_logic_vector(to_unsigned(213, 8)),
			3712 => std_logic_vector(to_unsigned(149, 8)),
			3713 => std_logic_vector(to_unsigned(121, 8)),
			3714 => std_logic_vector(to_unsigned(96, 8)),
			3715 => std_logic_vector(to_unsigned(178, 8)),
			3716 => std_logic_vector(to_unsigned(15, 8)),
			3717 => std_logic_vector(to_unsigned(65, 8)),
			3718 => std_logic_vector(to_unsigned(11, 8)),
			3719 => std_logic_vector(to_unsigned(118, 8)),
			3720 => std_logic_vector(to_unsigned(93, 8)),
			3721 => std_logic_vector(to_unsigned(205, 8)),
			3722 => std_logic_vector(to_unsigned(199, 8)),
			3723 => std_logic_vector(to_unsigned(84, 8)),
			3724 => std_logic_vector(to_unsigned(166, 8)),
			3725 => std_logic_vector(to_unsigned(118, 8)),
			3726 => std_logic_vector(to_unsigned(125, 8)),
			3727 => std_logic_vector(to_unsigned(228, 8)),
			3728 => std_logic_vector(to_unsigned(255, 8)),
			3729 => std_logic_vector(to_unsigned(251, 8)),
			3730 => std_logic_vector(to_unsigned(72, 8)),
			3731 => std_logic_vector(to_unsigned(153, 8)),
			3732 => std_logic_vector(to_unsigned(156, 8)),
			3733 => std_logic_vector(to_unsigned(146, 8)),
			3734 => std_logic_vector(to_unsigned(37, 8)),
			3735 => std_logic_vector(to_unsigned(231, 8)),
			3736 => std_logic_vector(to_unsigned(85, 8)),
			3737 => std_logic_vector(to_unsigned(176, 8)),
			3738 => std_logic_vector(to_unsigned(65, 8)),
			3739 => std_logic_vector(to_unsigned(115, 8)),
			3740 => std_logic_vector(to_unsigned(114, 8)),
			3741 => std_logic_vector(to_unsigned(235, 8)),
			3742 => std_logic_vector(to_unsigned(148, 8)),
			3743 => std_logic_vector(to_unsigned(68, 8)),
			3744 => std_logic_vector(to_unsigned(122, 8)),
			3745 => std_logic_vector(to_unsigned(59, 8)),
			3746 => std_logic_vector(to_unsigned(119, 8)),
			3747 => std_logic_vector(to_unsigned(49, 8)),
			3748 => std_logic_vector(to_unsigned(105, 8)),
			3749 => std_logic_vector(to_unsigned(100, 8)),
			3750 => std_logic_vector(to_unsigned(127, 8)),
			3751 => std_logic_vector(to_unsigned(23, 8)),
			3752 => std_logic_vector(to_unsigned(139, 8)),
			3753 => std_logic_vector(to_unsigned(232, 8)),
			3754 => std_logic_vector(to_unsigned(131, 8)),
			3755 => std_logic_vector(to_unsigned(243, 8)),
			3756 => std_logic_vector(to_unsigned(150, 8)),
			3757 => std_logic_vector(to_unsigned(16, 8)),
			3758 => std_logic_vector(to_unsigned(192, 8)),
			3759 => std_logic_vector(to_unsigned(107, 8)),
			3760 => std_logic_vector(to_unsigned(88, 8)),
			3761 => std_logic_vector(to_unsigned(61, 8)),
			3762 => std_logic_vector(to_unsigned(28, 8)),
			3763 => std_logic_vector(to_unsigned(166, 8)),
			3764 => std_logic_vector(to_unsigned(104, 8)),
			3765 => std_logic_vector(to_unsigned(250, 8)),
			3766 => std_logic_vector(to_unsigned(179, 8)),
			3767 => std_logic_vector(to_unsigned(59, 8)),
			3768 => std_logic_vector(to_unsigned(77, 8)),
			3769 => std_logic_vector(to_unsigned(169, 8)),
			3770 => std_logic_vector(to_unsigned(254, 8)),
			3771 => std_logic_vector(to_unsigned(138, 8)),
			3772 => std_logic_vector(to_unsigned(18, 8)),
			3773 => std_logic_vector(to_unsigned(3, 8)),
			3774 => std_logic_vector(to_unsigned(34, 8)),
			3775 => std_logic_vector(to_unsigned(55, 8)),
			3776 => std_logic_vector(to_unsigned(173, 8)),
			3777 => std_logic_vector(to_unsigned(144, 8)),
			3778 => std_logic_vector(to_unsigned(46, 8)),
			3779 => std_logic_vector(to_unsigned(97, 8)),
			3780 => std_logic_vector(to_unsigned(228, 8)),
			3781 => std_logic_vector(to_unsigned(187, 8)),
			3782 => std_logic_vector(to_unsigned(151, 8)),
			3783 => std_logic_vector(to_unsigned(224, 8)),
			3784 => std_logic_vector(to_unsigned(236, 8)),
			3785 => std_logic_vector(to_unsigned(96, 8)),
			3786 => std_logic_vector(to_unsigned(153, 8)),
			3787 => std_logic_vector(to_unsigned(188, 8)),
			3788 => std_logic_vector(to_unsigned(2, 8)),
			3789 => std_logic_vector(to_unsigned(147, 8)),
			3790 => std_logic_vector(to_unsigned(203, 8)),
			3791 => std_logic_vector(to_unsigned(50, 8)),
			3792 => std_logic_vector(to_unsigned(19, 8)),
			3793 => std_logic_vector(to_unsigned(146, 8)),
			3794 => std_logic_vector(to_unsigned(6, 8)),
			3795 => std_logic_vector(to_unsigned(50, 8)),
			3796 => std_logic_vector(to_unsigned(93, 8)),
			3797 => std_logic_vector(to_unsigned(123, 8)),
			3798 => std_logic_vector(to_unsigned(94, 8)),
			3799 => std_logic_vector(to_unsigned(115, 8)),
			3800 => std_logic_vector(to_unsigned(201, 8)),
			3801 => std_logic_vector(to_unsigned(176, 8)),
			3802 => std_logic_vector(to_unsigned(93, 8)),
			3803 => std_logic_vector(to_unsigned(48, 8)),
			3804 => std_logic_vector(to_unsigned(90, 8)),
			3805 => std_logic_vector(to_unsigned(180, 8)),
			3806 => std_logic_vector(to_unsigned(126, 8)),
			3807 => std_logic_vector(to_unsigned(245, 8)),
			3808 => std_logic_vector(to_unsigned(44, 8)),
			3809 => std_logic_vector(to_unsigned(191, 8)),
			3810 => std_logic_vector(to_unsigned(253, 8)),
			3811 => std_logic_vector(to_unsigned(26, 8)),
			3812 => std_logic_vector(to_unsigned(241, 8)),
			3813 => std_logic_vector(to_unsigned(3, 8)),
			3814 => std_logic_vector(to_unsigned(118, 8)),
			3815 => std_logic_vector(to_unsigned(170, 8)),
			3816 => std_logic_vector(to_unsigned(31, 8)),
			3817 => std_logic_vector(to_unsigned(133, 8)),
			3818 => std_logic_vector(to_unsigned(0, 8)),
			3819 => std_logic_vector(to_unsigned(237, 8)),
			3820 => std_logic_vector(to_unsigned(23, 8)),
			3821 => std_logic_vector(to_unsigned(41, 8)),
			3822 => std_logic_vector(to_unsigned(168, 8)),
			3823 => std_logic_vector(to_unsigned(135, 8)),
			3824 => std_logic_vector(to_unsigned(226, 8)),
			3825 => std_logic_vector(to_unsigned(72, 8)),
			3826 => std_logic_vector(to_unsigned(6, 8)),
			3827 => std_logic_vector(to_unsigned(52, 8)),
			3828 => std_logic_vector(to_unsigned(102, 8)),
			3829 => std_logic_vector(to_unsigned(93, 8)),
			3830 => std_logic_vector(to_unsigned(1, 8)),
			3831 => std_logic_vector(to_unsigned(106, 8)),
			3832 => std_logic_vector(to_unsigned(13, 8)),
			3833 => std_logic_vector(to_unsigned(2, 8)),
			3834 => std_logic_vector(to_unsigned(140, 8)),
			3835 => std_logic_vector(to_unsigned(148, 8)),
			3836 => std_logic_vector(to_unsigned(92, 8)),
			3837 => std_logic_vector(to_unsigned(188, 8)),
			3838 => std_logic_vector(to_unsigned(168, 8)),
			3839 => std_logic_vector(to_unsigned(147, 8)),
			3840 => std_logic_vector(to_unsigned(36, 8)),
			3841 => std_logic_vector(to_unsigned(74, 8)),
			3842 => std_logic_vector(to_unsigned(9, 8)),
			3843 => std_logic_vector(to_unsigned(109, 8)),
			3844 => std_logic_vector(to_unsigned(195, 8)),
			3845 => std_logic_vector(to_unsigned(69, 8)),
			3846 => std_logic_vector(to_unsigned(222, 8)),
			3847 => std_logic_vector(to_unsigned(68, 8)),
			3848 => std_logic_vector(to_unsigned(179, 8)),
			3849 => std_logic_vector(to_unsigned(35, 8)),
			3850 => std_logic_vector(to_unsigned(36, 8)),
			3851 => std_logic_vector(to_unsigned(250, 8)),
			3852 => std_logic_vector(to_unsigned(219, 8)),
			3853 => std_logic_vector(to_unsigned(41, 8)),
			3854 => std_logic_vector(to_unsigned(185, 8)),
			3855 => std_logic_vector(to_unsigned(153, 8)),
			3856 => std_logic_vector(to_unsigned(5, 8)),
			3857 => std_logic_vector(to_unsigned(145, 8)),
			3858 => std_logic_vector(to_unsigned(103, 8)),
			3859 => std_logic_vector(to_unsigned(2, 8)),
			3860 => std_logic_vector(to_unsigned(33, 8)),
			3861 => std_logic_vector(to_unsigned(249, 8)),
			3862 => std_logic_vector(to_unsigned(254, 8)),
			3863 => std_logic_vector(to_unsigned(172, 8)),
			3864 => std_logic_vector(to_unsigned(89, 8)),
			3865 => std_logic_vector(to_unsigned(139, 8)),
			3866 => std_logic_vector(to_unsigned(185, 8)),
			3867 => std_logic_vector(to_unsigned(69, 8)),
			3868 => std_logic_vector(to_unsigned(130, 8)),
			3869 => std_logic_vector(to_unsigned(216, 8)),
			3870 => std_logic_vector(to_unsigned(200, 8)),
			3871 => std_logic_vector(to_unsigned(113, 8)),
			3872 => std_logic_vector(to_unsigned(169, 8)),
			3873 => std_logic_vector(to_unsigned(81, 8)),
			3874 => std_logic_vector(to_unsigned(213, 8)),
			3875 => std_logic_vector(to_unsigned(135, 8)),
			3876 => std_logic_vector(to_unsigned(47, 8)),
			3877 => std_logic_vector(to_unsigned(23, 8)),
			3878 => std_logic_vector(to_unsigned(35, 8)),
			3879 => std_logic_vector(to_unsigned(146, 8)),
			3880 => std_logic_vector(to_unsigned(191, 8)),
			3881 => std_logic_vector(to_unsigned(211, 8)),
			3882 => std_logic_vector(to_unsigned(214, 8)),
			3883 => std_logic_vector(to_unsigned(71, 8)),
			3884 => std_logic_vector(to_unsigned(77, 8)),
			3885 => std_logic_vector(to_unsigned(226, 8)),
			3886 => std_logic_vector(to_unsigned(144, 8)),
			3887 => std_logic_vector(to_unsigned(243, 8)),
			3888 => std_logic_vector(to_unsigned(213, 8)),
			3889 => std_logic_vector(to_unsigned(146, 8)),
			3890 => std_logic_vector(to_unsigned(168, 8)),
			3891 => std_logic_vector(to_unsigned(126, 8)),
			3892 => std_logic_vector(to_unsigned(231, 8)),
			3893 => std_logic_vector(to_unsigned(205, 8)),
			3894 => std_logic_vector(to_unsigned(81, 8)),
			3895 => std_logic_vector(to_unsigned(7, 8)),
			3896 => std_logic_vector(to_unsigned(96, 8)),
			3897 => std_logic_vector(to_unsigned(250, 8)),
			3898 => std_logic_vector(to_unsigned(53, 8)),
			3899 => std_logic_vector(to_unsigned(64, 8)),
			3900 => std_logic_vector(to_unsigned(207, 8)),
			3901 => std_logic_vector(to_unsigned(184, 8)),
			3902 => std_logic_vector(to_unsigned(126, 8)),
			3903 => std_logic_vector(to_unsigned(10, 8)),
			3904 => std_logic_vector(to_unsigned(40, 8)),
			3905 => std_logic_vector(to_unsigned(216, 8)),
			3906 => std_logic_vector(to_unsigned(147, 8)),
			3907 => std_logic_vector(to_unsigned(180, 8)),
			3908 => std_logic_vector(to_unsigned(80, 8)),
			3909 => std_logic_vector(to_unsigned(139, 8)),
			3910 => std_logic_vector(to_unsigned(47, 8)),
			3911 => std_logic_vector(to_unsigned(182, 8)),
			3912 => std_logic_vector(to_unsigned(15, 8)),
			3913 => std_logic_vector(to_unsigned(207, 8)),
			3914 => std_logic_vector(to_unsigned(169, 8)),
			3915 => std_logic_vector(to_unsigned(180, 8)),
			3916 => std_logic_vector(to_unsigned(158, 8)),
			3917 => std_logic_vector(to_unsigned(169, 8)),
			3918 => std_logic_vector(to_unsigned(185, 8)),
			3919 => std_logic_vector(to_unsigned(195, 8)),
			3920 => std_logic_vector(to_unsigned(86, 8)),
			3921 => std_logic_vector(to_unsigned(153, 8)),
			3922 => std_logic_vector(to_unsigned(105, 8)),
			3923 => std_logic_vector(to_unsigned(154, 8)),
			3924 => std_logic_vector(to_unsigned(36, 8)),
			3925 => std_logic_vector(to_unsigned(241, 8)),
			3926 => std_logic_vector(to_unsigned(10, 8)),
			3927 => std_logic_vector(to_unsigned(178, 8)),
			3928 => std_logic_vector(to_unsigned(221, 8)),
			3929 => std_logic_vector(to_unsigned(26, 8)),
			3930 => std_logic_vector(to_unsigned(108, 8)),
			3931 => std_logic_vector(to_unsigned(179, 8)),
			3932 => std_logic_vector(to_unsigned(229, 8)),
			3933 => std_logic_vector(to_unsigned(154, 8)),
			3934 => std_logic_vector(to_unsigned(95, 8)),
			3935 => std_logic_vector(to_unsigned(228, 8)),
			3936 => std_logic_vector(to_unsigned(170, 8)),
			3937 => std_logic_vector(to_unsigned(5, 8)),
			3938 => std_logic_vector(to_unsigned(173, 8)),
			3939 => std_logic_vector(to_unsigned(11, 8)),
			3940 => std_logic_vector(to_unsigned(155, 8)),
			3941 => std_logic_vector(to_unsigned(169, 8)),
			3942 => std_logic_vector(to_unsigned(135, 8)),
			3943 => std_logic_vector(to_unsigned(127, 8)),
			3944 => std_logic_vector(to_unsigned(233, 8)),
			3945 => std_logic_vector(to_unsigned(96, 8)),
			3946 => std_logic_vector(to_unsigned(119, 8)),
			3947 => std_logic_vector(to_unsigned(91, 8)),
			3948 => std_logic_vector(to_unsigned(43, 8)),
			3949 => std_logic_vector(to_unsigned(163, 8)),
			3950 => std_logic_vector(to_unsigned(7, 8)),
			3951 => std_logic_vector(to_unsigned(127, 8)),
			3952 => std_logic_vector(to_unsigned(30, 8)),
			3953 => std_logic_vector(to_unsigned(241, 8)),
			3954 => std_logic_vector(to_unsigned(211, 8)),
			3955 => std_logic_vector(to_unsigned(167, 8)),
			3956 => std_logic_vector(to_unsigned(9, 8)),
			3957 => std_logic_vector(to_unsigned(250, 8)),
			3958 => std_logic_vector(to_unsigned(236, 8)),
			3959 => std_logic_vector(to_unsigned(249, 8)),
			3960 => std_logic_vector(to_unsigned(123, 8)),
			3961 => std_logic_vector(to_unsigned(81, 8)),
			3962 => std_logic_vector(to_unsigned(245, 8)),
			3963 => std_logic_vector(to_unsigned(31, 8)),
			3964 => std_logic_vector(to_unsigned(130, 8)),
			3965 => std_logic_vector(to_unsigned(62, 8)),
			3966 => std_logic_vector(to_unsigned(18, 8)),
			3967 => std_logic_vector(to_unsigned(241, 8)),
			3968 => std_logic_vector(to_unsigned(44, 8)),
			3969 => std_logic_vector(to_unsigned(147, 8)),
			3970 => std_logic_vector(to_unsigned(230, 8)),
			3971 => std_logic_vector(to_unsigned(25, 8)),
			3972 => std_logic_vector(to_unsigned(121, 8)),
			3973 => std_logic_vector(to_unsigned(73, 8)),
			3974 => std_logic_vector(to_unsigned(247, 8)),
			3975 => std_logic_vector(to_unsigned(217, 8)),
			3976 => std_logic_vector(to_unsigned(108, 8)),
			3977 => std_logic_vector(to_unsigned(10, 8)),
			3978 => std_logic_vector(to_unsigned(10, 8)),
			3979 => std_logic_vector(to_unsigned(65, 8)),
			3980 => std_logic_vector(to_unsigned(14, 8)),
			3981 => std_logic_vector(to_unsigned(115, 8)),
			3982 => std_logic_vector(to_unsigned(248, 8)),
			3983 => std_logic_vector(to_unsigned(147, 8)),
			3984 => std_logic_vector(to_unsigned(155, 8)),
			3985 => std_logic_vector(to_unsigned(71, 8)),
			3986 => std_logic_vector(to_unsigned(91, 8)),
			3987 => std_logic_vector(to_unsigned(2, 8)),
			3988 => std_logic_vector(to_unsigned(222, 8)),
			3989 => std_logic_vector(to_unsigned(68, 8)),
			3990 => std_logic_vector(to_unsigned(25, 8)),
			3991 => std_logic_vector(to_unsigned(43, 8)),
			3992 => std_logic_vector(to_unsigned(142, 8)),
			3993 => std_logic_vector(to_unsigned(229, 8)),
			3994 => std_logic_vector(to_unsigned(23, 8)),
			3995 => std_logic_vector(to_unsigned(226, 8)),
			3996 => std_logic_vector(to_unsigned(238, 8)),
			3997 => std_logic_vector(to_unsigned(28, 8)),
			3998 => std_logic_vector(to_unsigned(53, 8)),
			3999 => std_logic_vector(to_unsigned(178, 8)),
			4000 => std_logic_vector(to_unsigned(72, 8)),
			4001 => std_logic_vector(to_unsigned(3, 8)),
			4002 => std_logic_vector(to_unsigned(248, 8)),
			4003 => std_logic_vector(to_unsigned(123, 8)),
			4004 => std_logic_vector(to_unsigned(252, 8)),
			4005 => std_logic_vector(to_unsigned(18, 8)),
			4006 => std_logic_vector(to_unsigned(164, 8)),
			4007 => std_logic_vector(to_unsigned(173, 8)),
			4008 => std_logic_vector(to_unsigned(162, 8)),
			4009 => std_logic_vector(to_unsigned(158, 8)),
			4010 => std_logic_vector(to_unsigned(83, 8)),
			4011 => std_logic_vector(to_unsigned(128, 8)),
			4012 => std_logic_vector(to_unsigned(236, 8)),
			4013 => std_logic_vector(to_unsigned(88, 8)),
			4014 => std_logic_vector(to_unsigned(189, 8)),
			4015 => std_logic_vector(to_unsigned(220, 8)),
			4016 => std_logic_vector(to_unsigned(109, 8)),
			4017 => std_logic_vector(to_unsigned(66, 8)),
			4018 => std_logic_vector(to_unsigned(39, 8)),
			4019 => std_logic_vector(to_unsigned(52, 8)),
			4020 => std_logic_vector(to_unsigned(148, 8)),
			4021 => std_logic_vector(to_unsigned(101, 8)),
			4022 => std_logic_vector(to_unsigned(106, 8)),
			4023 => std_logic_vector(to_unsigned(101, 8)),
			4024 => std_logic_vector(to_unsigned(200, 8)),
			4025 => std_logic_vector(to_unsigned(40, 8)),
			4026 => std_logic_vector(to_unsigned(32, 8)),
			4027 => std_logic_vector(to_unsigned(65, 8)),
			4028 => std_logic_vector(to_unsigned(146, 8)),
			4029 => std_logic_vector(to_unsigned(17, 8)),
			4030 => std_logic_vector(to_unsigned(218, 8)),
			4031 => std_logic_vector(to_unsigned(167, 8)),
			4032 => std_logic_vector(to_unsigned(91, 8)),
			4033 => std_logic_vector(to_unsigned(196, 8)),
			4034 => std_logic_vector(to_unsigned(249, 8)),
			4035 => std_logic_vector(to_unsigned(188, 8)),
			4036 => std_logic_vector(to_unsigned(4, 8)),
			4037 => std_logic_vector(to_unsigned(151, 8)),
			4038 => std_logic_vector(to_unsigned(20, 8)),
			4039 => std_logic_vector(to_unsigned(129, 8)),
			4040 => std_logic_vector(to_unsigned(57, 8)),
			4041 => std_logic_vector(to_unsigned(1, 8)),
			4042 => std_logic_vector(to_unsigned(121, 8)),
			4043 => std_logic_vector(to_unsigned(167, 8)),
			4044 => std_logic_vector(to_unsigned(240, 8)),
			4045 => std_logic_vector(to_unsigned(210, 8)),
			4046 => std_logic_vector(to_unsigned(18, 8)),
			4047 => std_logic_vector(to_unsigned(34, 8)),
			4048 => std_logic_vector(to_unsigned(87, 8)),
			4049 => std_logic_vector(to_unsigned(49, 8)),
			4050 => std_logic_vector(to_unsigned(101, 8)),
			4051 => std_logic_vector(to_unsigned(141, 8)),
			4052 => std_logic_vector(to_unsigned(95, 8)),
			4053 => std_logic_vector(to_unsigned(111, 8)),
			4054 => std_logic_vector(to_unsigned(253, 8)),
			4055 => std_logic_vector(to_unsigned(253, 8)),
			4056 => std_logic_vector(to_unsigned(125, 8)),
			4057 => std_logic_vector(to_unsigned(137, 8)),
			4058 => std_logic_vector(to_unsigned(102, 8)),
			4059 => std_logic_vector(to_unsigned(222, 8)),
			4060 => std_logic_vector(to_unsigned(136, 8)),
			4061 => std_logic_vector(to_unsigned(254, 8)),
			4062 => std_logic_vector(to_unsigned(71, 8)),
			4063 => std_logic_vector(to_unsigned(122, 8)),
			4064 => std_logic_vector(to_unsigned(236, 8)),
			4065 => std_logic_vector(to_unsigned(235, 8)),
			4066 => std_logic_vector(to_unsigned(51, 8)),
			4067 => std_logic_vector(to_unsigned(56, 8)),
			4068 => std_logic_vector(to_unsigned(205, 8)),
			4069 => std_logic_vector(to_unsigned(216, 8)),
			4070 => std_logic_vector(to_unsigned(22, 8)),
			4071 => std_logic_vector(to_unsigned(210, 8)),
			4072 => std_logic_vector(to_unsigned(60, 8)),
			4073 => std_logic_vector(to_unsigned(55, 8)),
			4074 => std_logic_vector(to_unsigned(142, 8)),
			4075 => std_logic_vector(to_unsigned(70, 8)),
			4076 => std_logic_vector(to_unsigned(108, 8)),
			4077 => std_logic_vector(to_unsigned(230, 8)),
			4078 => std_logic_vector(to_unsigned(140, 8)),
			4079 => std_logic_vector(to_unsigned(145, 8)),
			4080 => std_logic_vector(to_unsigned(61, 8)),
			4081 => std_logic_vector(to_unsigned(98, 8)),
			4082 => std_logic_vector(to_unsigned(5, 8)),
			4083 => std_logic_vector(to_unsigned(124, 8)),
			4084 => std_logic_vector(to_unsigned(37, 8)),
			4085 => std_logic_vector(to_unsigned(62, 8)),
			4086 => std_logic_vector(to_unsigned(102, 8)),
			4087 => std_logic_vector(to_unsigned(205, 8)),
			4088 => std_logic_vector(to_unsigned(5, 8)),
			4089 => std_logic_vector(to_unsigned(45, 8)),
			4090 => std_logic_vector(to_unsigned(215, 8)),
			4091 => std_logic_vector(to_unsigned(151, 8)),
			4092 => std_logic_vector(to_unsigned(119, 8)),
			4093 => std_logic_vector(to_unsigned(171, 8)),
			4094 => std_logic_vector(to_unsigned(126, 8)),
			4095 => std_logic_vector(to_unsigned(73, 8)),
			4096 => std_logic_vector(to_unsigned(163, 8)),
			4097 => std_logic_vector(to_unsigned(3, 8)),
			4098 => std_logic_vector(to_unsigned(120, 8)),
			4099 => std_logic_vector(to_unsigned(100, 8)),
			4100 => std_logic_vector(to_unsigned(149, 8)),
			4101 => std_logic_vector(to_unsigned(92, 8)),
			4102 => std_logic_vector(to_unsigned(227, 8)),
			4103 => std_logic_vector(to_unsigned(219, 8)),
			4104 => std_logic_vector(to_unsigned(81, 8)),
			4105 => std_logic_vector(to_unsigned(16, 8)),
			4106 => std_logic_vector(to_unsigned(169, 8)),
			4107 => std_logic_vector(to_unsigned(194, 8)),
			4108 => std_logic_vector(to_unsigned(161, 8)),
			4109 => std_logic_vector(to_unsigned(3, 8)),
			4110 => std_logic_vector(to_unsigned(149, 8)),
			4111 => std_logic_vector(to_unsigned(42, 8)),
			4112 => std_logic_vector(to_unsigned(164, 8)),
			4113 => std_logic_vector(to_unsigned(24, 8)),
			4114 => std_logic_vector(to_unsigned(19, 8)),
			4115 => std_logic_vector(to_unsigned(253, 8)),
			4116 => std_logic_vector(to_unsigned(144, 8)),
			4117 => std_logic_vector(to_unsigned(236, 8)),
			4118 => std_logic_vector(to_unsigned(47, 8)),
			4119 => std_logic_vector(to_unsigned(186, 8)),
			4120 => std_logic_vector(to_unsigned(168, 8)),
			4121 => std_logic_vector(to_unsigned(73, 8)),
			4122 => std_logic_vector(to_unsigned(74, 8)),
			4123 => std_logic_vector(to_unsigned(92, 8)),
			4124 => std_logic_vector(to_unsigned(242, 8)),
			4125 => std_logic_vector(to_unsigned(250, 8)),
			4126 => std_logic_vector(to_unsigned(200, 8)),
			4127 => std_logic_vector(to_unsigned(201, 8)),
			4128 => std_logic_vector(to_unsigned(88, 8)),
			4129 => std_logic_vector(to_unsigned(121, 8)),
			4130 => std_logic_vector(to_unsigned(83, 8)),
			4131 => std_logic_vector(to_unsigned(115, 8)),
			4132 => std_logic_vector(to_unsigned(75, 8)),
			4133 => std_logic_vector(to_unsigned(122, 8)),
			4134 => std_logic_vector(to_unsigned(124, 8)),
			4135 => std_logic_vector(to_unsigned(224, 8)),
			4136 => std_logic_vector(to_unsigned(245, 8)),
			4137 => std_logic_vector(to_unsigned(183, 8)),
			4138 => std_logic_vector(to_unsigned(70, 8)),
			4139 => std_logic_vector(to_unsigned(212, 8)),
			4140 => std_logic_vector(to_unsigned(77, 8)),
			4141 => std_logic_vector(to_unsigned(159, 8)),
			4142 => std_logic_vector(to_unsigned(55, 8)),
			4143 => std_logic_vector(to_unsigned(68, 8)),
			4144 => std_logic_vector(to_unsigned(12, 8)),
			4145 => std_logic_vector(to_unsigned(252, 8)),
			4146 => std_logic_vector(to_unsigned(135, 8)),
			4147 => std_logic_vector(to_unsigned(52, 8)),
			4148 => std_logic_vector(to_unsigned(148, 8)),
			4149 => std_logic_vector(to_unsigned(207, 8)),
			4150 => std_logic_vector(to_unsigned(54, 8)),
			4151 => std_logic_vector(to_unsigned(247, 8)),
			4152 => std_logic_vector(to_unsigned(33, 8)),
			4153 => std_logic_vector(to_unsigned(153, 8)),
			4154 => std_logic_vector(to_unsigned(155, 8)),
			4155 => std_logic_vector(to_unsigned(20, 8)),
			4156 => std_logic_vector(to_unsigned(242, 8)),
			4157 => std_logic_vector(to_unsigned(14, 8)),
			4158 => std_logic_vector(to_unsigned(44, 8)),
			4159 => std_logic_vector(to_unsigned(75, 8)),
			4160 => std_logic_vector(to_unsigned(94, 8)),
			4161 => std_logic_vector(to_unsigned(169, 8)),
			4162 => std_logic_vector(to_unsigned(64, 8)),
			4163 => std_logic_vector(to_unsigned(232, 8)),
			4164 => std_logic_vector(to_unsigned(128, 8)),
			4165 => std_logic_vector(to_unsigned(24, 8)),
			4166 => std_logic_vector(to_unsigned(200, 8)),
			4167 => std_logic_vector(to_unsigned(211, 8)),
			4168 => std_logic_vector(to_unsigned(199, 8)),
			4169 => std_logic_vector(to_unsigned(63, 8)),
			4170 => std_logic_vector(to_unsigned(66, 8)),
			4171 => std_logic_vector(to_unsigned(75, 8)),
			4172 => std_logic_vector(to_unsigned(5, 8)),
			4173 => std_logic_vector(to_unsigned(146, 8)),
			4174 => std_logic_vector(to_unsigned(58, 8)),
			4175 => std_logic_vector(to_unsigned(45, 8)),
			4176 => std_logic_vector(to_unsigned(18, 8)),
			4177 => std_logic_vector(to_unsigned(171, 8)),
			4178 => std_logic_vector(to_unsigned(226, 8)),
			4179 => std_logic_vector(to_unsigned(168, 8)),
			4180 => std_logic_vector(to_unsigned(62, 8)),
			4181 => std_logic_vector(to_unsigned(41, 8)),
			4182 => std_logic_vector(to_unsigned(133, 8)),
			4183 => std_logic_vector(to_unsigned(93, 8)),
			4184 => std_logic_vector(to_unsigned(79, 8)),
			4185 => std_logic_vector(to_unsigned(147, 8)),
			4186 => std_logic_vector(to_unsigned(87, 8)),
			4187 => std_logic_vector(to_unsigned(170, 8)),
			4188 => std_logic_vector(to_unsigned(95, 8)),
			4189 => std_logic_vector(to_unsigned(165, 8)),
			4190 => std_logic_vector(to_unsigned(191, 8)),
			4191 => std_logic_vector(to_unsigned(106, 8)),
			4192 => std_logic_vector(to_unsigned(176, 8)),
			4193 => std_logic_vector(to_unsigned(163, 8)),
			4194 => std_logic_vector(to_unsigned(30, 8)),
			4195 => std_logic_vector(to_unsigned(31, 8)),
			4196 => std_logic_vector(to_unsigned(88, 8)),
			4197 => std_logic_vector(to_unsigned(85, 8)),
			4198 => std_logic_vector(to_unsigned(55, 8)),
			4199 => std_logic_vector(to_unsigned(155, 8)),
			4200 => std_logic_vector(to_unsigned(227, 8)),
			4201 => std_logic_vector(to_unsigned(204, 8)),
			4202 => std_logic_vector(to_unsigned(99, 8)),
			4203 => std_logic_vector(to_unsigned(228, 8)),
			4204 => std_logic_vector(to_unsigned(4, 8)),
			4205 => std_logic_vector(to_unsigned(145, 8)),
			4206 => std_logic_vector(to_unsigned(93, 8)),
			4207 => std_logic_vector(to_unsigned(213, 8)),
			4208 => std_logic_vector(to_unsigned(57, 8)),
			4209 => std_logic_vector(to_unsigned(244, 8)),
			4210 => std_logic_vector(to_unsigned(162, 8)),
			4211 => std_logic_vector(to_unsigned(179, 8)),
			4212 => std_logic_vector(to_unsigned(214, 8)),
			4213 => std_logic_vector(to_unsigned(17, 8)),
			4214 => std_logic_vector(to_unsigned(154, 8)),
			4215 => std_logic_vector(to_unsigned(236, 8)),
			4216 => std_logic_vector(to_unsigned(157, 8)),
			4217 => std_logic_vector(to_unsigned(85, 8)),
			4218 => std_logic_vector(to_unsigned(168, 8)),
			4219 => std_logic_vector(to_unsigned(74, 8)),
			4220 => std_logic_vector(to_unsigned(197, 8)),
			4221 => std_logic_vector(to_unsigned(50, 8)),
			4222 => std_logic_vector(to_unsigned(111, 8)),
			4223 => std_logic_vector(to_unsigned(133, 8)),
			4224 => std_logic_vector(to_unsigned(39, 8)),
			4225 => std_logic_vector(to_unsigned(251, 8)),
			4226 => std_logic_vector(to_unsigned(230, 8)),
			4227 => std_logic_vector(to_unsigned(141, 8)),
			4228 => std_logic_vector(to_unsigned(67, 8)),
			4229 => std_logic_vector(to_unsigned(64, 8)),
			4230 => std_logic_vector(to_unsigned(0, 8)),
			4231 => std_logic_vector(to_unsigned(77, 8)),
			4232 => std_logic_vector(to_unsigned(212, 8)),
			4233 => std_logic_vector(to_unsigned(73, 8)),
			4234 => std_logic_vector(to_unsigned(15, 8)),
			4235 => std_logic_vector(to_unsigned(240, 8)),
			4236 => std_logic_vector(to_unsigned(29, 8)),
			4237 => std_logic_vector(to_unsigned(218, 8)),
			4238 => std_logic_vector(to_unsigned(50, 8)),
			4239 => std_logic_vector(to_unsigned(8, 8)),
			4240 => std_logic_vector(to_unsigned(255, 8)),
			4241 => std_logic_vector(to_unsigned(93, 8)),
			4242 => std_logic_vector(to_unsigned(83, 8)),
			4243 => std_logic_vector(to_unsigned(253, 8)),
			4244 => std_logic_vector(to_unsigned(65, 8)),
			4245 => std_logic_vector(to_unsigned(182, 8)),
			4246 => std_logic_vector(to_unsigned(224, 8)),
			4247 => std_logic_vector(to_unsigned(24, 8)),
			4248 => std_logic_vector(to_unsigned(237, 8)),
			4249 => std_logic_vector(to_unsigned(208, 8)),
			4250 => std_logic_vector(to_unsigned(236, 8)),
			4251 => std_logic_vector(to_unsigned(24, 8)),
			4252 => std_logic_vector(to_unsigned(202, 8)),
			4253 => std_logic_vector(to_unsigned(189, 8)),
			4254 => std_logic_vector(to_unsigned(157, 8)),
			4255 => std_logic_vector(to_unsigned(77, 8)),
			4256 => std_logic_vector(to_unsigned(174, 8)),
			4257 => std_logic_vector(to_unsigned(241, 8)),
			4258 => std_logic_vector(to_unsigned(247, 8)),
			4259 => std_logic_vector(to_unsigned(245, 8)),
			4260 => std_logic_vector(to_unsigned(43, 8)),
			4261 => std_logic_vector(to_unsigned(145, 8)),
			4262 => std_logic_vector(to_unsigned(247, 8)),
			4263 => std_logic_vector(to_unsigned(233, 8)),
			4264 => std_logic_vector(to_unsigned(78, 8)),
			4265 => std_logic_vector(to_unsigned(111, 8)),
			4266 => std_logic_vector(to_unsigned(75, 8)),
			4267 => std_logic_vector(to_unsigned(228, 8)),
			4268 => std_logic_vector(to_unsigned(255, 8)),
			4269 => std_logic_vector(to_unsigned(187, 8)),
			4270 => std_logic_vector(to_unsigned(201, 8)),
			4271 => std_logic_vector(to_unsigned(219, 8)),
			4272 => std_logic_vector(to_unsigned(49, 8)),
			4273 => std_logic_vector(to_unsigned(179, 8)),
			4274 => std_logic_vector(to_unsigned(138, 8)),
			4275 => std_logic_vector(to_unsigned(99, 8)),
			4276 => std_logic_vector(to_unsigned(76, 8)),
			4277 => std_logic_vector(to_unsigned(224, 8)),
			4278 => std_logic_vector(to_unsigned(107, 8)),
			4279 => std_logic_vector(to_unsigned(80, 8)),
			4280 => std_logic_vector(to_unsigned(245, 8)),
			4281 => std_logic_vector(to_unsigned(172, 8)),
			4282 => std_logic_vector(to_unsigned(182, 8)),
			4283 => std_logic_vector(to_unsigned(154, 8)),
			4284 => std_logic_vector(to_unsigned(23, 8)),
			4285 => std_logic_vector(to_unsigned(208, 8)),
			4286 => std_logic_vector(to_unsigned(210, 8)),
			4287 => std_logic_vector(to_unsigned(235, 8)),
			4288 => std_logic_vector(to_unsigned(155, 8)),
			4289 => std_logic_vector(to_unsigned(57, 8)),
			4290 => std_logic_vector(to_unsigned(189, 8)),
			4291 => std_logic_vector(to_unsigned(254, 8)),
			4292 => std_logic_vector(to_unsigned(122, 8)),
			4293 => std_logic_vector(to_unsigned(215, 8)),
			4294 => std_logic_vector(to_unsigned(34, 8)),
			4295 => std_logic_vector(to_unsigned(188, 8)),
			4296 => std_logic_vector(to_unsigned(118, 8)),
			4297 => std_logic_vector(to_unsigned(39, 8)),
			4298 => std_logic_vector(to_unsigned(59, 8)),
			4299 => std_logic_vector(to_unsigned(205, 8)),
			4300 => std_logic_vector(to_unsigned(50, 8)),
			4301 => std_logic_vector(to_unsigned(101, 8)),
			4302 => std_logic_vector(to_unsigned(106, 8)),
			4303 => std_logic_vector(to_unsigned(7, 8)),
			4304 => std_logic_vector(to_unsigned(196, 8)),
			4305 => std_logic_vector(to_unsigned(226, 8)),
			4306 => std_logic_vector(to_unsigned(56, 8)),
			4307 => std_logic_vector(to_unsigned(102, 8)),
			4308 => std_logic_vector(to_unsigned(57, 8)),
			4309 => std_logic_vector(to_unsigned(81, 8)),
			4310 => std_logic_vector(to_unsigned(220, 8)),
			4311 => std_logic_vector(to_unsigned(209, 8)),
			4312 => std_logic_vector(to_unsigned(171, 8)),
			4313 => std_logic_vector(to_unsigned(192, 8)),
			4314 => std_logic_vector(to_unsigned(184, 8)),
			4315 => std_logic_vector(to_unsigned(128, 8)),
			4316 => std_logic_vector(to_unsigned(126, 8)),
			4317 => std_logic_vector(to_unsigned(12, 8)),
			4318 => std_logic_vector(to_unsigned(2, 8)),
			4319 => std_logic_vector(to_unsigned(56, 8)),
			4320 => std_logic_vector(to_unsigned(12, 8)),
			4321 => std_logic_vector(to_unsigned(236, 8)),
			4322 => std_logic_vector(to_unsigned(144, 8)),
			4323 => std_logic_vector(to_unsigned(138, 8)),
			4324 => std_logic_vector(to_unsigned(216, 8)),
			4325 => std_logic_vector(to_unsigned(105, 8)),
			4326 => std_logic_vector(to_unsigned(85, 8)),
			4327 => std_logic_vector(to_unsigned(148, 8)),
			4328 => std_logic_vector(to_unsigned(179, 8)),
			4329 => std_logic_vector(to_unsigned(125, 8)),
			4330 => std_logic_vector(to_unsigned(6, 8)),
			4331 => std_logic_vector(to_unsigned(142, 8)),
			4332 => std_logic_vector(to_unsigned(34, 8)),
			4333 => std_logic_vector(to_unsigned(231, 8)),
			4334 => std_logic_vector(to_unsigned(76, 8)),
			4335 => std_logic_vector(to_unsigned(128, 8)),
			4336 => std_logic_vector(to_unsigned(217, 8)),
			4337 => std_logic_vector(to_unsigned(225, 8)),
			4338 => std_logic_vector(to_unsigned(208, 8)),
			4339 => std_logic_vector(to_unsigned(123, 8)),
			4340 => std_logic_vector(to_unsigned(153, 8)),
			4341 => std_logic_vector(to_unsigned(160, 8)),
			4342 => std_logic_vector(to_unsigned(117, 8)),
			4343 => std_logic_vector(to_unsigned(250, 8)),
			4344 => std_logic_vector(to_unsigned(83, 8)),
			4345 => std_logic_vector(to_unsigned(157, 8)),
			4346 => std_logic_vector(to_unsigned(243, 8)),
			4347 => std_logic_vector(to_unsigned(251, 8)),
			4348 => std_logic_vector(to_unsigned(63, 8)),
			4349 => std_logic_vector(to_unsigned(78, 8)),
			4350 => std_logic_vector(to_unsigned(84, 8)),
			4351 => std_logic_vector(to_unsigned(171, 8)),
			4352 => std_logic_vector(to_unsigned(57, 8)),
			4353 => std_logic_vector(to_unsigned(119, 8)),
			4354 => std_logic_vector(to_unsigned(221, 8)),
			4355 => std_logic_vector(to_unsigned(9, 8)),
			4356 => std_logic_vector(to_unsigned(86, 8)),
			4357 => std_logic_vector(to_unsigned(55, 8)),
			4358 => std_logic_vector(to_unsigned(117, 8)),
			4359 => std_logic_vector(to_unsigned(93, 8)),
			4360 => std_logic_vector(to_unsigned(16, 8)),
			4361 => std_logic_vector(to_unsigned(235, 8)),
			4362 => std_logic_vector(to_unsigned(24, 8)),
			4363 => std_logic_vector(to_unsigned(93, 8)),
			4364 => std_logic_vector(to_unsigned(108, 8)),
			4365 => std_logic_vector(to_unsigned(165, 8)),
			4366 => std_logic_vector(to_unsigned(169, 8)),
			4367 => std_logic_vector(to_unsigned(61, 8)),
			4368 => std_logic_vector(to_unsigned(4, 8)),
			4369 => std_logic_vector(to_unsigned(88, 8)),
			4370 => std_logic_vector(to_unsigned(204, 8)),
			4371 => std_logic_vector(to_unsigned(181, 8)),
			4372 => std_logic_vector(to_unsigned(61, 8)),
			4373 => std_logic_vector(to_unsigned(50, 8)),
			4374 => std_logic_vector(to_unsigned(71, 8)),
			4375 => std_logic_vector(to_unsigned(80, 8)),
			4376 => std_logic_vector(to_unsigned(207, 8)),
			4377 => std_logic_vector(to_unsigned(194, 8)),
			4378 => std_logic_vector(to_unsigned(40, 8)),
			4379 => std_logic_vector(to_unsigned(56, 8)),
			4380 => std_logic_vector(to_unsigned(11, 8)),
			4381 => std_logic_vector(to_unsigned(26, 8)),
			4382 => std_logic_vector(to_unsigned(219, 8)),
			4383 => std_logic_vector(to_unsigned(87, 8)),
			4384 => std_logic_vector(to_unsigned(207, 8)),
			4385 => std_logic_vector(to_unsigned(98, 8)),
			4386 => std_logic_vector(to_unsigned(19, 8)),
			4387 => std_logic_vector(to_unsigned(158, 8)),
			4388 => std_logic_vector(to_unsigned(9, 8)),
			4389 => std_logic_vector(to_unsigned(251, 8)),
			4390 => std_logic_vector(to_unsigned(132, 8)),
			4391 => std_logic_vector(to_unsigned(123, 8)),
			4392 => std_logic_vector(to_unsigned(73, 8)),
			4393 => std_logic_vector(to_unsigned(23, 8)),
			4394 => std_logic_vector(to_unsigned(44, 8)),
			4395 => std_logic_vector(to_unsigned(99, 8)),
			4396 => std_logic_vector(to_unsigned(65, 8)),
			4397 => std_logic_vector(to_unsigned(231, 8)),
			4398 => std_logic_vector(to_unsigned(218, 8)),
			4399 => std_logic_vector(to_unsigned(184, 8)),
			4400 => std_logic_vector(to_unsigned(76, 8)),
			4401 => std_logic_vector(to_unsigned(187, 8)),
			4402 => std_logic_vector(to_unsigned(88, 8)),
			4403 => std_logic_vector(to_unsigned(206, 8)),
			4404 => std_logic_vector(to_unsigned(6, 8)),
			4405 => std_logic_vector(to_unsigned(175, 8)),
			4406 => std_logic_vector(to_unsigned(74, 8)),
			4407 => std_logic_vector(to_unsigned(110, 8)),
			4408 => std_logic_vector(to_unsigned(56, 8)),
			4409 => std_logic_vector(to_unsigned(161, 8)),
			4410 => std_logic_vector(to_unsigned(183, 8)),
			4411 => std_logic_vector(to_unsigned(206, 8)),
			4412 => std_logic_vector(to_unsigned(83, 8)),
			4413 => std_logic_vector(to_unsigned(248, 8)),
			4414 => std_logic_vector(to_unsigned(73, 8)),
			4415 => std_logic_vector(to_unsigned(106, 8)),
			4416 => std_logic_vector(to_unsigned(47, 8)),
			4417 => std_logic_vector(to_unsigned(95, 8)),
			4418 => std_logic_vector(to_unsigned(170, 8)),
			4419 => std_logic_vector(to_unsigned(222, 8)),
			4420 => std_logic_vector(to_unsigned(11, 8)),
			4421 => std_logic_vector(to_unsigned(242, 8)),
			4422 => std_logic_vector(to_unsigned(76, 8)),
			4423 => std_logic_vector(to_unsigned(66, 8)),
			4424 => std_logic_vector(to_unsigned(174, 8)),
			4425 => std_logic_vector(to_unsigned(171, 8)),
			4426 => std_logic_vector(to_unsigned(46, 8)),
			4427 => std_logic_vector(to_unsigned(23, 8)),
			4428 => std_logic_vector(to_unsigned(150, 8)),
			4429 => std_logic_vector(to_unsigned(199, 8)),
			4430 => std_logic_vector(to_unsigned(253, 8)),
			4431 => std_logic_vector(to_unsigned(142, 8)),
			4432 => std_logic_vector(to_unsigned(251, 8)),
			4433 => std_logic_vector(to_unsigned(12, 8)),
			4434 => std_logic_vector(to_unsigned(49, 8)),
			4435 => std_logic_vector(to_unsigned(94, 8)),
			4436 => std_logic_vector(to_unsigned(130, 8)),
			4437 => std_logic_vector(to_unsigned(230, 8)),
			4438 => std_logic_vector(to_unsigned(229, 8)),
			4439 => std_logic_vector(to_unsigned(178, 8)),
			4440 => std_logic_vector(to_unsigned(14, 8)),
			4441 => std_logic_vector(to_unsigned(32, 8)),
			4442 => std_logic_vector(to_unsigned(150, 8)),
			4443 => std_logic_vector(to_unsigned(71, 8)),
			4444 => std_logic_vector(to_unsigned(208, 8)),
			4445 => std_logic_vector(to_unsigned(199, 8)),
			4446 => std_logic_vector(to_unsigned(124, 8)),
			4447 => std_logic_vector(to_unsigned(71, 8)),
			4448 => std_logic_vector(to_unsigned(203, 8)),
			4449 => std_logic_vector(to_unsigned(127, 8)),
			4450 => std_logic_vector(to_unsigned(99, 8)),
			4451 => std_logic_vector(to_unsigned(111, 8)),
			4452 => std_logic_vector(to_unsigned(48, 8)),
			4453 => std_logic_vector(to_unsigned(112, 8)),
			4454 => std_logic_vector(to_unsigned(75, 8)),
			4455 => std_logic_vector(to_unsigned(44, 8)),
			4456 => std_logic_vector(to_unsigned(174, 8)),
			4457 => std_logic_vector(to_unsigned(71, 8)),
			4458 => std_logic_vector(to_unsigned(90, 8)),
			4459 => std_logic_vector(to_unsigned(131, 8)),
			4460 => std_logic_vector(to_unsigned(204, 8)),
			4461 => std_logic_vector(to_unsigned(209, 8)),
			4462 => std_logic_vector(to_unsigned(234, 8)),
			4463 => std_logic_vector(to_unsigned(49, 8)),
			4464 => std_logic_vector(to_unsigned(255, 8)),
			4465 => std_logic_vector(to_unsigned(148, 8)),
			4466 => std_logic_vector(to_unsigned(50, 8)),
			4467 => std_logic_vector(to_unsigned(247, 8)),
			4468 => std_logic_vector(to_unsigned(203, 8)),
			4469 => std_logic_vector(to_unsigned(221, 8)),
			4470 => std_logic_vector(to_unsigned(187, 8)),
			4471 => std_logic_vector(to_unsigned(199, 8)),
			4472 => std_logic_vector(to_unsigned(213, 8)),
			4473 => std_logic_vector(to_unsigned(92, 8)),
			4474 => std_logic_vector(to_unsigned(160, 8)),
			4475 => std_logic_vector(to_unsigned(44, 8)),
			4476 => std_logic_vector(to_unsigned(165, 8)),
			4477 => std_logic_vector(to_unsigned(38, 8)),
			4478 => std_logic_vector(to_unsigned(68, 8)),
			4479 => std_logic_vector(to_unsigned(36, 8)),
			4480 => std_logic_vector(to_unsigned(84, 8)),
			4481 => std_logic_vector(to_unsigned(161, 8)),
			4482 => std_logic_vector(to_unsigned(23, 8)),
			4483 => std_logic_vector(to_unsigned(111, 8)),
			4484 => std_logic_vector(to_unsigned(137, 8)),
			4485 => std_logic_vector(to_unsigned(87, 8)),
			4486 => std_logic_vector(to_unsigned(41, 8)),
			4487 => std_logic_vector(to_unsigned(24, 8)),
			4488 => std_logic_vector(to_unsigned(222, 8)),
			4489 => std_logic_vector(to_unsigned(28, 8)),
			4490 => std_logic_vector(to_unsigned(111, 8)),
			4491 => std_logic_vector(to_unsigned(71, 8)),
			4492 => std_logic_vector(to_unsigned(221, 8)),
			4493 => std_logic_vector(to_unsigned(41, 8)),
			4494 => std_logic_vector(to_unsigned(178, 8)),
			4495 => std_logic_vector(to_unsigned(242, 8)),
			4496 => std_logic_vector(to_unsigned(38, 8)),
			4497 => std_logic_vector(to_unsigned(144, 8)),
			4498 => std_logic_vector(to_unsigned(60, 8)),
			4499 => std_logic_vector(to_unsigned(165, 8)),
			4500 => std_logic_vector(to_unsigned(125, 8)),
			4501 => std_logic_vector(to_unsigned(10, 8)),
			4502 => std_logic_vector(to_unsigned(99, 8)),
			4503 => std_logic_vector(to_unsigned(19, 8)),
			4504 => std_logic_vector(to_unsigned(148, 8)),
			4505 => std_logic_vector(to_unsigned(253, 8)),
			4506 => std_logic_vector(to_unsigned(29, 8)),
			4507 => std_logic_vector(to_unsigned(238, 8)),
			4508 => std_logic_vector(to_unsigned(20, 8)),
			4509 => std_logic_vector(to_unsigned(217, 8)),
			4510 => std_logic_vector(to_unsigned(157, 8)),
			4511 => std_logic_vector(to_unsigned(86, 8)),
			4512 => std_logic_vector(to_unsigned(229, 8)),
			4513 => std_logic_vector(to_unsigned(59, 8)),
			4514 => std_logic_vector(to_unsigned(125, 8)),
			4515 => std_logic_vector(to_unsigned(227, 8)),
			4516 => std_logic_vector(to_unsigned(139, 8)),
			4517 => std_logic_vector(to_unsigned(131, 8)),
			4518 => std_logic_vector(to_unsigned(219, 8)),
			4519 => std_logic_vector(to_unsigned(104, 8)),
			4520 => std_logic_vector(to_unsigned(203, 8)),
			4521 => std_logic_vector(to_unsigned(0, 8)),
			4522 => std_logic_vector(to_unsigned(179, 8)),
			4523 => std_logic_vector(to_unsigned(254, 8)),
			4524 => std_logic_vector(to_unsigned(132, 8)),
			4525 => std_logic_vector(to_unsigned(9, 8)),
			4526 => std_logic_vector(to_unsigned(239, 8)),
			4527 => std_logic_vector(to_unsigned(120, 8)),
			4528 => std_logic_vector(to_unsigned(23, 8)),
			4529 => std_logic_vector(to_unsigned(86, 8)),
			4530 => std_logic_vector(to_unsigned(94, 8)),
			4531 => std_logic_vector(to_unsigned(212, 8)),
			4532 => std_logic_vector(to_unsigned(12, 8)),
			4533 => std_logic_vector(to_unsigned(242, 8)),
			4534 => std_logic_vector(to_unsigned(5, 8)),
			4535 => std_logic_vector(to_unsigned(17, 8)),
			4536 => std_logic_vector(to_unsigned(83, 8)),
			4537 => std_logic_vector(to_unsigned(50, 8)),
			4538 => std_logic_vector(to_unsigned(106, 8)),
			4539 => std_logic_vector(to_unsigned(0, 8)),
			4540 => std_logic_vector(to_unsigned(145, 8)),
			4541 => std_logic_vector(to_unsigned(166, 8)),
			4542 => std_logic_vector(to_unsigned(31, 8)),
			4543 => std_logic_vector(to_unsigned(161, 8)),
			4544 => std_logic_vector(to_unsigned(61, 8)),
			4545 => std_logic_vector(to_unsigned(56, 8)),
			4546 => std_logic_vector(to_unsigned(232, 8)),
			4547 => std_logic_vector(to_unsigned(212, 8)),
			4548 => std_logic_vector(to_unsigned(76, 8)),
			4549 => std_logic_vector(to_unsigned(50, 8)),
			4550 => std_logic_vector(to_unsigned(136, 8)),
			4551 => std_logic_vector(to_unsigned(137, 8)),
			4552 => std_logic_vector(to_unsigned(253, 8)),
			4553 => std_logic_vector(to_unsigned(70, 8)),
			4554 => std_logic_vector(to_unsigned(202, 8)),
			4555 => std_logic_vector(to_unsigned(97, 8)),
			4556 => std_logic_vector(to_unsigned(94, 8)),
			4557 => std_logic_vector(to_unsigned(3, 8)),
			4558 => std_logic_vector(to_unsigned(48, 8)),
			4559 => std_logic_vector(to_unsigned(86, 8)),
			4560 => std_logic_vector(to_unsigned(231, 8)),
			4561 => std_logic_vector(to_unsigned(63, 8)),
			4562 => std_logic_vector(to_unsigned(41, 8)),
			4563 => std_logic_vector(to_unsigned(15, 8)),
			4564 => std_logic_vector(to_unsigned(81, 8)),
			4565 => std_logic_vector(to_unsigned(162, 8)),
			4566 => std_logic_vector(to_unsigned(62, 8)),
			4567 => std_logic_vector(to_unsigned(37, 8)),
			4568 => std_logic_vector(to_unsigned(87, 8)),
			4569 => std_logic_vector(to_unsigned(41, 8)),
			4570 => std_logic_vector(to_unsigned(115, 8)),
			4571 => std_logic_vector(to_unsigned(99, 8)),
			4572 => std_logic_vector(to_unsigned(87, 8)),
			4573 => std_logic_vector(to_unsigned(91, 8)),
			4574 => std_logic_vector(to_unsigned(217, 8)),
			4575 => std_logic_vector(to_unsigned(141, 8)),
			4576 => std_logic_vector(to_unsigned(156, 8)),
			4577 => std_logic_vector(to_unsigned(173, 8)),
			4578 => std_logic_vector(to_unsigned(158, 8)),
			4579 => std_logic_vector(to_unsigned(8, 8)),
			4580 => std_logic_vector(to_unsigned(187, 8)),
			4581 => std_logic_vector(to_unsigned(250, 8)),
			4582 => std_logic_vector(to_unsigned(176, 8)),
			4583 => std_logic_vector(to_unsigned(105, 8)),
			4584 => std_logic_vector(to_unsigned(223, 8)),
			4585 => std_logic_vector(to_unsigned(247, 8)),
			4586 => std_logic_vector(to_unsigned(79, 8)),
			4587 => std_logic_vector(to_unsigned(71, 8)),
			4588 => std_logic_vector(to_unsigned(167, 8)),
			4589 => std_logic_vector(to_unsigned(11, 8)),
			4590 => std_logic_vector(to_unsigned(28, 8)),
			4591 => std_logic_vector(to_unsigned(137, 8)),
			4592 => std_logic_vector(to_unsigned(90, 8)),
			4593 => std_logic_vector(to_unsigned(91, 8)),
			4594 => std_logic_vector(to_unsigned(18, 8)),
			4595 => std_logic_vector(to_unsigned(127, 8)),
			4596 => std_logic_vector(to_unsigned(129, 8)),
			4597 => std_logic_vector(to_unsigned(24, 8)),
			4598 => std_logic_vector(to_unsigned(231, 8)),
			4599 => std_logic_vector(to_unsigned(94, 8)),
			4600 => std_logic_vector(to_unsigned(235, 8)),
			4601 => std_logic_vector(to_unsigned(159, 8)),
			4602 => std_logic_vector(to_unsigned(168, 8)),
			4603 => std_logic_vector(to_unsigned(175, 8)),
			4604 => std_logic_vector(to_unsigned(8, 8)),
			4605 => std_logic_vector(to_unsigned(234, 8)),
			4606 => std_logic_vector(to_unsigned(41, 8)),
			4607 => std_logic_vector(to_unsigned(236, 8)),
			4608 => std_logic_vector(to_unsigned(237, 8)),
			4609 => std_logic_vector(to_unsigned(97, 8)),
			4610 => std_logic_vector(to_unsigned(199, 8)),
			4611 => std_logic_vector(to_unsigned(166, 8)),
			4612 => std_logic_vector(to_unsigned(209, 8)),
			4613 => std_logic_vector(to_unsigned(189, 8)),
			4614 => std_logic_vector(to_unsigned(149, 8)),
			4615 => std_logic_vector(to_unsigned(151, 8)),
			4616 => std_logic_vector(to_unsigned(162, 8)),
			4617 => std_logic_vector(to_unsigned(9, 8)),
			4618 => std_logic_vector(to_unsigned(162, 8)),
			4619 => std_logic_vector(to_unsigned(9, 8)),
			4620 => std_logic_vector(to_unsigned(129, 8)),
			4621 => std_logic_vector(to_unsigned(114, 8)),
			4622 => std_logic_vector(to_unsigned(15, 8)),
			4623 => std_logic_vector(to_unsigned(196, 8)),
			4624 => std_logic_vector(to_unsigned(193, 8)),
			4625 => std_logic_vector(to_unsigned(119, 8)),
			4626 => std_logic_vector(to_unsigned(169, 8)),
			4627 => std_logic_vector(to_unsigned(170, 8)),
			4628 => std_logic_vector(to_unsigned(39, 8)),
			4629 => std_logic_vector(to_unsigned(253, 8)),
			4630 => std_logic_vector(to_unsigned(7, 8)),
			4631 => std_logic_vector(to_unsigned(175, 8)),
			4632 => std_logic_vector(to_unsigned(233, 8)),
			4633 => std_logic_vector(to_unsigned(140, 8)),
			4634 => std_logic_vector(to_unsigned(81, 8)),
			4635 => std_logic_vector(to_unsigned(191, 8)),
			4636 => std_logic_vector(to_unsigned(25, 8)),
			4637 => std_logic_vector(to_unsigned(95, 8)),
			4638 => std_logic_vector(to_unsigned(71, 8)),
			4639 => std_logic_vector(to_unsigned(172, 8)),
			4640 => std_logic_vector(to_unsigned(154, 8)),
			4641 => std_logic_vector(to_unsigned(6, 8)),
			4642 => std_logic_vector(to_unsigned(220, 8)),
			4643 => std_logic_vector(to_unsigned(96, 8)),
			4644 => std_logic_vector(to_unsigned(83, 8)),
			4645 => std_logic_vector(to_unsigned(153, 8)),
			4646 => std_logic_vector(to_unsigned(228, 8)),
			4647 => std_logic_vector(to_unsigned(20, 8)),
			4648 => std_logic_vector(to_unsigned(120, 8)),
			4649 => std_logic_vector(to_unsigned(159, 8)),
			4650 => std_logic_vector(to_unsigned(142, 8)),
			4651 => std_logic_vector(to_unsigned(172, 8)),
			4652 => std_logic_vector(to_unsigned(3, 8)),
			4653 => std_logic_vector(to_unsigned(166, 8)),
			4654 => std_logic_vector(to_unsigned(0, 8)),
			4655 => std_logic_vector(to_unsigned(89, 8)),
			4656 => std_logic_vector(to_unsigned(105, 8)),
			4657 => std_logic_vector(to_unsigned(72, 8)),
			4658 => std_logic_vector(to_unsigned(92, 8)),
			4659 => std_logic_vector(to_unsigned(81, 8)),
			4660 => std_logic_vector(to_unsigned(206, 8)),
			4661 => std_logic_vector(to_unsigned(179, 8)),
			4662 => std_logic_vector(to_unsigned(14, 8)),
			4663 => std_logic_vector(to_unsigned(28, 8)),
			4664 => std_logic_vector(to_unsigned(102, 8)),
			4665 => std_logic_vector(to_unsigned(189, 8)),
			4666 => std_logic_vector(to_unsigned(157, 8)),
			4667 => std_logic_vector(to_unsigned(202, 8)),
			4668 => std_logic_vector(to_unsigned(111, 8)),
			4669 => std_logic_vector(to_unsigned(121, 8)),
			4670 => std_logic_vector(to_unsigned(209, 8)),
			4671 => std_logic_vector(to_unsigned(11, 8)),
			4672 => std_logic_vector(to_unsigned(127, 8)),
			4673 => std_logic_vector(to_unsigned(148, 8)),
			4674 => std_logic_vector(to_unsigned(184, 8)),
			4675 => std_logic_vector(to_unsigned(16, 8)),
			4676 => std_logic_vector(to_unsigned(139, 8)),
			4677 => std_logic_vector(to_unsigned(186, 8)),
			4678 => std_logic_vector(to_unsigned(242, 8)),
			4679 => std_logic_vector(to_unsigned(237, 8)),
			4680 => std_logic_vector(to_unsigned(150, 8)),
			4681 => std_logic_vector(to_unsigned(253, 8)),
			4682 => std_logic_vector(to_unsigned(170, 8)),
			4683 => std_logic_vector(to_unsigned(120, 8)),
			4684 => std_logic_vector(to_unsigned(108, 8)),
			4685 => std_logic_vector(to_unsigned(19, 8)),
			4686 => std_logic_vector(to_unsigned(137, 8)),
			4687 => std_logic_vector(to_unsigned(152, 8)),
			4688 => std_logic_vector(to_unsigned(74, 8)),
			4689 => std_logic_vector(to_unsigned(130, 8)),
			4690 => std_logic_vector(to_unsigned(119, 8)),
			4691 => std_logic_vector(to_unsigned(150, 8)),
			4692 => std_logic_vector(to_unsigned(107, 8)),
			4693 => std_logic_vector(to_unsigned(25, 8)),
			4694 => std_logic_vector(to_unsigned(3, 8)),
			4695 => std_logic_vector(to_unsigned(108, 8)),
			4696 => std_logic_vector(to_unsigned(41, 8)),
			4697 => std_logic_vector(to_unsigned(42, 8)),
			4698 => std_logic_vector(to_unsigned(171, 8)),
			4699 => std_logic_vector(to_unsigned(170, 8)),
			4700 => std_logic_vector(to_unsigned(190, 8)),
			4701 => std_logic_vector(to_unsigned(168, 8)),
			4702 => std_logic_vector(to_unsigned(156, 8)),
			4703 => std_logic_vector(to_unsigned(203, 8)),
			4704 => std_logic_vector(to_unsigned(252, 8)),
			4705 => std_logic_vector(to_unsigned(167, 8)),
			4706 => std_logic_vector(to_unsigned(104, 8)),
			4707 => std_logic_vector(to_unsigned(119, 8)),
			4708 => std_logic_vector(to_unsigned(240, 8)),
			4709 => std_logic_vector(to_unsigned(82, 8)),
			4710 => std_logic_vector(to_unsigned(230, 8)),
			4711 => std_logic_vector(to_unsigned(240, 8)),
			4712 => std_logic_vector(to_unsigned(161, 8)),
			4713 => std_logic_vector(to_unsigned(140, 8)),
			4714 => std_logic_vector(to_unsigned(201, 8)),
			4715 => std_logic_vector(to_unsigned(80, 8)),
			4716 => std_logic_vector(to_unsigned(142, 8)),
			4717 => std_logic_vector(to_unsigned(211, 8)),
			4718 => std_logic_vector(to_unsigned(109, 8)),
			4719 => std_logic_vector(to_unsigned(232, 8)),
			4720 => std_logic_vector(to_unsigned(183, 8)),
			4721 => std_logic_vector(to_unsigned(88, 8)),
			4722 => std_logic_vector(to_unsigned(38, 8)),
			4723 => std_logic_vector(to_unsigned(73, 8)),
			4724 => std_logic_vector(to_unsigned(217, 8)),
			4725 => std_logic_vector(to_unsigned(103, 8)),
			4726 => std_logic_vector(to_unsigned(158, 8)),
			4727 => std_logic_vector(to_unsigned(209, 8)),
			4728 => std_logic_vector(to_unsigned(93, 8)),
			4729 => std_logic_vector(to_unsigned(253, 8)),
			4730 => std_logic_vector(to_unsigned(227, 8)),
			4731 => std_logic_vector(to_unsigned(173, 8)),
			4732 => std_logic_vector(to_unsigned(108, 8)),
			4733 => std_logic_vector(to_unsigned(94, 8)),
			4734 => std_logic_vector(to_unsigned(195, 8)),
			4735 => std_logic_vector(to_unsigned(232, 8)),
			4736 => std_logic_vector(to_unsigned(114, 8)),
			4737 => std_logic_vector(to_unsigned(114, 8)),
			4738 => std_logic_vector(to_unsigned(176, 8)),
			4739 => std_logic_vector(to_unsigned(191, 8)),
			4740 => std_logic_vector(to_unsigned(76, 8)),
			4741 => std_logic_vector(to_unsigned(215, 8)),
			4742 => std_logic_vector(to_unsigned(215, 8)),
			4743 => std_logic_vector(to_unsigned(150, 8)),
			4744 => std_logic_vector(to_unsigned(51, 8)),
			4745 => std_logic_vector(to_unsigned(99, 8)),
			4746 => std_logic_vector(to_unsigned(233, 8)),
			4747 => std_logic_vector(to_unsigned(217, 8)),
			4748 => std_logic_vector(to_unsigned(27, 8)),
			4749 => std_logic_vector(to_unsigned(193, 8)),
			4750 => std_logic_vector(to_unsigned(49, 8)),
			4751 => std_logic_vector(to_unsigned(63, 8)),
			4752 => std_logic_vector(to_unsigned(78, 8)),
			4753 => std_logic_vector(to_unsigned(148, 8)),
			4754 => std_logic_vector(to_unsigned(22, 8)),
			4755 => std_logic_vector(to_unsigned(97, 8)),
			4756 => std_logic_vector(to_unsigned(237, 8)),
			4757 => std_logic_vector(to_unsigned(30, 8)),
			4758 => std_logic_vector(to_unsigned(225, 8)),
			4759 => std_logic_vector(to_unsigned(235, 8)),
			4760 => std_logic_vector(to_unsigned(34, 8)),
			4761 => std_logic_vector(to_unsigned(220, 8)),
			4762 => std_logic_vector(to_unsigned(45, 8)),
			4763 => std_logic_vector(to_unsigned(103, 8)),
			4764 => std_logic_vector(to_unsigned(2, 8)),
			4765 => std_logic_vector(to_unsigned(154, 8)),
			4766 => std_logic_vector(to_unsigned(123, 8)),
			4767 => std_logic_vector(to_unsigned(149, 8)),
			4768 => std_logic_vector(to_unsigned(73, 8)),
			4769 => std_logic_vector(to_unsigned(199, 8)),
			4770 => std_logic_vector(to_unsigned(172, 8)),
			4771 => std_logic_vector(to_unsigned(142, 8)),
			4772 => std_logic_vector(to_unsigned(112, 8)),
			4773 => std_logic_vector(to_unsigned(92, 8)),
			4774 => std_logic_vector(to_unsigned(207, 8)),
			4775 => std_logic_vector(to_unsigned(238, 8)),
			4776 => std_logic_vector(to_unsigned(17, 8)),
			4777 => std_logic_vector(to_unsigned(122, 8)),
			4778 => std_logic_vector(to_unsigned(48, 8)),
			4779 => std_logic_vector(to_unsigned(87, 8)),
			4780 => std_logic_vector(to_unsigned(74, 8)),
			4781 => std_logic_vector(to_unsigned(90, 8)),
			4782 => std_logic_vector(to_unsigned(181, 8)),
			4783 => std_logic_vector(to_unsigned(183, 8)),
			4784 => std_logic_vector(to_unsigned(57, 8)),
			4785 => std_logic_vector(to_unsigned(234, 8)),
			4786 => std_logic_vector(to_unsigned(227, 8)),
			4787 => std_logic_vector(to_unsigned(201, 8)),
			4788 => std_logic_vector(to_unsigned(249, 8)),
			4789 => std_logic_vector(to_unsigned(244, 8)),
			4790 => std_logic_vector(to_unsigned(50, 8)),
			4791 => std_logic_vector(to_unsigned(6, 8)),
			4792 => std_logic_vector(to_unsigned(94, 8)),
			4793 => std_logic_vector(to_unsigned(249, 8)),
			4794 => std_logic_vector(to_unsigned(169, 8)),
			4795 => std_logic_vector(to_unsigned(160, 8)),
			4796 => std_logic_vector(to_unsigned(74, 8)),
			4797 => std_logic_vector(to_unsigned(85, 8)),
			4798 => std_logic_vector(to_unsigned(125, 8)),
			4799 => std_logic_vector(to_unsigned(193, 8)),
			4800 => std_logic_vector(to_unsigned(81, 8)),
			4801 => std_logic_vector(to_unsigned(212, 8)),
			4802 => std_logic_vector(to_unsigned(99, 8)),
			4803 => std_logic_vector(to_unsigned(176, 8)),
			4804 => std_logic_vector(to_unsigned(174, 8)),
			4805 => std_logic_vector(to_unsigned(133, 8)),
			4806 => std_logic_vector(to_unsigned(180, 8)),
			4807 => std_logic_vector(to_unsigned(116, 8)),
			4808 => std_logic_vector(to_unsigned(219, 8)),
			4809 => std_logic_vector(to_unsigned(71, 8)),
			4810 => std_logic_vector(to_unsigned(18, 8)),
			4811 => std_logic_vector(to_unsigned(192, 8)),
			4812 => std_logic_vector(to_unsigned(137, 8)),
			4813 => std_logic_vector(to_unsigned(26, 8)),
			4814 => std_logic_vector(to_unsigned(49, 8)),
			4815 => std_logic_vector(to_unsigned(204, 8)),
			4816 => std_logic_vector(to_unsigned(43, 8)),
			4817 => std_logic_vector(to_unsigned(134, 8)),
			4818 => std_logic_vector(to_unsigned(210, 8)),
			4819 => std_logic_vector(to_unsigned(141, 8)),
			4820 => std_logic_vector(to_unsigned(215, 8)),
			4821 => std_logic_vector(to_unsigned(172, 8)),
			4822 => std_logic_vector(to_unsigned(48, 8)),
			4823 => std_logic_vector(to_unsigned(231, 8)),
			4824 => std_logic_vector(to_unsigned(179, 8)),
			4825 => std_logic_vector(to_unsigned(182, 8)),
			4826 => std_logic_vector(to_unsigned(56, 8)),
			4827 => std_logic_vector(to_unsigned(105, 8)),
			4828 => std_logic_vector(to_unsigned(95, 8)),
			4829 => std_logic_vector(to_unsigned(72, 8)),
			4830 => std_logic_vector(to_unsigned(136, 8)),
			4831 => std_logic_vector(to_unsigned(215, 8)),
			4832 => std_logic_vector(to_unsigned(81, 8)),
			4833 => std_logic_vector(to_unsigned(221, 8)),
			4834 => std_logic_vector(to_unsigned(66, 8)),
			4835 => std_logic_vector(to_unsigned(46, 8)),
			4836 => std_logic_vector(to_unsigned(116, 8)),
			4837 => std_logic_vector(to_unsigned(16, 8)),
			4838 => std_logic_vector(to_unsigned(97, 8)),
			4839 => std_logic_vector(to_unsigned(154, 8)),
			4840 => std_logic_vector(to_unsigned(95, 8)),
			4841 => std_logic_vector(to_unsigned(74, 8)),
			4842 => std_logic_vector(to_unsigned(86, 8)),
			4843 => std_logic_vector(to_unsigned(53, 8)),
			4844 => std_logic_vector(to_unsigned(20, 8)),
			4845 => std_logic_vector(to_unsigned(45, 8)),
			4846 => std_logic_vector(to_unsigned(113, 8)),
			4847 => std_logic_vector(to_unsigned(19, 8)),
			4848 => std_logic_vector(to_unsigned(242, 8)),
			4849 => std_logic_vector(to_unsigned(173, 8)),
			4850 => std_logic_vector(to_unsigned(233, 8)),
			4851 => std_logic_vector(to_unsigned(65, 8)),
			4852 => std_logic_vector(to_unsigned(152, 8)),
			4853 => std_logic_vector(to_unsigned(45, 8)),
			4854 => std_logic_vector(to_unsigned(172, 8)),
			4855 => std_logic_vector(to_unsigned(189, 8)),
			4856 => std_logic_vector(to_unsigned(129, 8)),
			4857 => std_logic_vector(to_unsigned(217, 8)),
			4858 => std_logic_vector(to_unsigned(119, 8)),
			4859 => std_logic_vector(to_unsigned(76, 8)),
			4860 => std_logic_vector(to_unsigned(87, 8)),
			4861 => std_logic_vector(to_unsigned(213, 8)),
			4862 => std_logic_vector(to_unsigned(61, 8)),
			4863 => std_logic_vector(to_unsigned(239, 8)),
			4864 => std_logic_vector(to_unsigned(220, 8)),
			4865 => std_logic_vector(to_unsigned(13, 8)),
			4866 => std_logic_vector(to_unsigned(190, 8)),
			4867 => std_logic_vector(to_unsigned(164, 8)),
			4868 => std_logic_vector(to_unsigned(93, 8)),
			4869 => std_logic_vector(to_unsigned(222, 8)),
			4870 => std_logic_vector(to_unsigned(91, 8)),
			4871 => std_logic_vector(to_unsigned(226, 8)),
			4872 => std_logic_vector(to_unsigned(39, 8)),
			4873 => std_logic_vector(to_unsigned(60, 8)),
			4874 => std_logic_vector(to_unsigned(122, 8)),
			4875 => std_logic_vector(to_unsigned(139, 8)),
			4876 => std_logic_vector(to_unsigned(141, 8)),
			4877 => std_logic_vector(to_unsigned(177, 8)),
			4878 => std_logic_vector(to_unsigned(16, 8)),
			4879 => std_logic_vector(to_unsigned(27, 8)),
			4880 => std_logic_vector(to_unsigned(88, 8)),
			4881 => std_logic_vector(to_unsigned(113, 8)),
			4882 => std_logic_vector(to_unsigned(98, 8)),
			4883 => std_logic_vector(to_unsigned(119, 8)),
			4884 => std_logic_vector(to_unsigned(252, 8)),
			4885 => std_logic_vector(to_unsigned(107, 8)),
			4886 => std_logic_vector(to_unsigned(241, 8)),
			4887 => std_logic_vector(to_unsigned(202, 8)),
			4888 => std_logic_vector(to_unsigned(199, 8)),
			4889 => std_logic_vector(to_unsigned(155, 8)),
			4890 => std_logic_vector(to_unsigned(7, 8)),
			4891 => std_logic_vector(to_unsigned(160, 8)),
			4892 => std_logic_vector(to_unsigned(30, 8)),
			4893 => std_logic_vector(to_unsigned(64, 8)),
			4894 => std_logic_vector(to_unsigned(117, 8)),
			4895 => std_logic_vector(to_unsigned(130, 8)),
			4896 => std_logic_vector(to_unsigned(61, 8)),
			4897 => std_logic_vector(to_unsigned(243, 8)),
			4898 => std_logic_vector(to_unsigned(96, 8)),
			4899 => std_logic_vector(to_unsigned(96, 8)),
			4900 => std_logic_vector(to_unsigned(103, 8)),
			4901 => std_logic_vector(to_unsigned(235, 8)),
			4902 => std_logic_vector(to_unsigned(41, 8)),
			4903 => std_logic_vector(to_unsigned(122, 8)),
			4904 => std_logic_vector(to_unsigned(190, 8)),
			4905 => std_logic_vector(to_unsigned(250, 8)),
			4906 => std_logic_vector(to_unsigned(164, 8)),
			4907 => std_logic_vector(to_unsigned(234, 8)),
			4908 => std_logic_vector(to_unsigned(125, 8)),
			4909 => std_logic_vector(to_unsigned(26, 8)),
			4910 => std_logic_vector(to_unsigned(243, 8)),
			4911 => std_logic_vector(to_unsigned(199, 8)),
			4912 => std_logic_vector(to_unsigned(253, 8)),
			4913 => std_logic_vector(to_unsigned(142, 8)),
			4914 => std_logic_vector(to_unsigned(171, 8)),
			4915 => std_logic_vector(to_unsigned(204, 8)),
			4916 => std_logic_vector(to_unsigned(124, 8)),
			4917 => std_logic_vector(to_unsigned(19, 8)),
			4918 => std_logic_vector(to_unsigned(34, 8)),
			4919 => std_logic_vector(to_unsigned(35, 8)),
			4920 => std_logic_vector(to_unsigned(10, 8)),
			4921 => std_logic_vector(to_unsigned(59, 8)),
			4922 => std_logic_vector(to_unsigned(39, 8)),
			4923 => std_logic_vector(to_unsigned(169, 8)),
			4924 => std_logic_vector(to_unsigned(180, 8)),
			4925 => std_logic_vector(to_unsigned(250, 8)),
			4926 => std_logic_vector(to_unsigned(142, 8)),
			4927 => std_logic_vector(to_unsigned(248, 8)),
			4928 => std_logic_vector(to_unsigned(67, 8)),
			4929 => std_logic_vector(to_unsigned(9, 8)),
			4930 => std_logic_vector(to_unsigned(105, 8)),
			4931 => std_logic_vector(to_unsigned(205, 8)),
			4932 => std_logic_vector(to_unsigned(10, 8)),
			4933 => std_logic_vector(to_unsigned(141, 8)),
			4934 => std_logic_vector(to_unsigned(135, 8)),
			4935 => std_logic_vector(to_unsigned(103, 8)),
			4936 => std_logic_vector(to_unsigned(230, 8)),
			4937 => std_logic_vector(to_unsigned(192, 8)),
			4938 => std_logic_vector(to_unsigned(48, 8)),
			4939 => std_logic_vector(to_unsigned(35, 8)),
			4940 => std_logic_vector(to_unsigned(114, 8)),
			4941 => std_logic_vector(to_unsigned(143, 8)),
			4942 => std_logic_vector(to_unsigned(101, 8)),
			4943 => std_logic_vector(to_unsigned(28, 8)),
			4944 => std_logic_vector(to_unsigned(168, 8)),
			4945 => std_logic_vector(to_unsigned(110, 8)),
			4946 => std_logic_vector(to_unsigned(27, 8)),
			4947 => std_logic_vector(to_unsigned(246, 8)),
			4948 => std_logic_vector(to_unsigned(219, 8)),
			4949 => std_logic_vector(to_unsigned(89, 8)),
			4950 => std_logic_vector(to_unsigned(136, 8)),
			4951 => std_logic_vector(to_unsigned(14, 8)),
			4952 => std_logic_vector(to_unsigned(143, 8)),
			4953 => std_logic_vector(to_unsigned(206, 8)),
			4954 => std_logic_vector(to_unsigned(215, 8)),
			4955 => std_logic_vector(to_unsigned(205, 8)),
			4956 => std_logic_vector(to_unsigned(71, 8)),
			4957 => std_logic_vector(to_unsigned(69, 8)),
			4958 => std_logic_vector(to_unsigned(134, 8)),
			4959 => std_logic_vector(to_unsigned(25, 8)),
			4960 => std_logic_vector(to_unsigned(84, 8)),
			4961 => std_logic_vector(to_unsigned(11, 8)),
			4962 => std_logic_vector(to_unsigned(50, 8)),
			4963 => std_logic_vector(to_unsigned(42, 8)),
			4964 => std_logic_vector(to_unsigned(179, 8)),
			4965 => std_logic_vector(to_unsigned(104, 8)),
			4966 => std_logic_vector(to_unsigned(231, 8)),
			4967 => std_logic_vector(to_unsigned(232, 8)),
			4968 => std_logic_vector(to_unsigned(71, 8)),
			4969 => std_logic_vector(to_unsigned(153, 8)),
			4970 => std_logic_vector(to_unsigned(101, 8)),
			4971 => std_logic_vector(to_unsigned(22, 8)),
			4972 => std_logic_vector(to_unsigned(145, 8)),
			4973 => std_logic_vector(to_unsigned(111, 8)),
			4974 => std_logic_vector(to_unsigned(44, 8)),
			4975 => std_logic_vector(to_unsigned(83, 8)),
			4976 => std_logic_vector(to_unsigned(254, 8)),
			4977 => std_logic_vector(to_unsigned(142, 8)),
			4978 => std_logic_vector(to_unsigned(143, 8)),
			4979 => std_logic_vector(to_unsigned(245, 8)),
			4980 => std_logic_vector(to_unsigned(231, 8)),
			4981 => std_logic_vector(to_unsigned(241, 8)),
			4982 => std_logic_vector(to_unsigned(195, 8)),
			4983 => std_logic_vector(to_unsigned(80, 8)),
			4984 => std_logic_vector(to_unsigned(53, 8)),
			4985 => std_logic_vector(to_unsigned(158, 8)),
			4986 => std_logic_vector(to_unsigned(88, 8)),
			4987 => std_logic_vector(to_unsigned(0, 8)),
			4988 => std_logic_vector(to_unsigned(229, 8)),
			4989 => std_logic_vector(to_unsigned(252, 8)),
			4990 => std_logic_vector(to_unsigned(217, 8)),
			4991 => std_logic_vector(to_unsigned(122, 8)),
			4992 => std_logic_vector(to_unsigned(173, 8)),
			4993 => std_logic_vector(to_unsigned(154, 8)),
			4994 => std_logic_vector(to_unsigned(219, 8)),
			4995 => std_logic_vector(to_unsigned(143, 8)),
			4996 => std_logic_vector(to_unsigned(87, 8)),
			4997 => std_logic_vector(to_unsigned(118, 8)),
			4998 => std_logic_vector(to_unsigned(182, 8)),
			4999 => std_logic_vector(to_unsigned(17, 8)),
			5000 => std_logic_vector(to_unsigned(165, 8)),
			5001 => std_logic_vector(to_unsigned(252, 8)),
			5002 => std_logic_vector(to_unsigned(189, 8)),
			5003 => std_logic_vector(to_unsigned(14, 8)),
			5004 => std_logic_vector(to_unsigned(55, 8)),
			5005 => std_logic_vector(to_unsigned(245, 8)),
			5006 => std_logic_vector(to_unsigned(205, 8)),
			5007 => std_logic_vector(to_unsigned(33, 8)),
			5008 => std_logic_vector(to_unsigned(97, 8)),
			5009 => std_logic_vector(to_unsigned(56, 8)),
			5010 => std_logic_vector(to_unsigned(183, 8)),
			5011 => std_logic_vector(to_unsigned(94, 8)),
			5012 => std_logic_vector(to_unsigned(94, 8)),
			5013 => std_logic_vector(to_unsigned(123, 8)),
			5014 => std_logic_vector(to_unsigned(20, 8)),
			5015 => std_logic_vector(to_unsigned(42, 8)),
			5016 => std_logic_vector(to_unsigned(71, 8)),
			5017 => std_logic_vector(to_unsigned(200, 8)),
			5018 => std_logic_vector(to_unsigned(2, 8)),
			5019 => std_logic_vector(to_unsigned(71, 8)),
			5020 => std_logic_vector(to_unsigned(225, 8)),
			5021 => std_logic_vector(to_unsigned(26, 8)),
			5022 => std_logic_vector(to_unsigned(186, 8)),
			5023 => std_logic_vector(to_unsigned(203, 8)),
			5024 => std_logic_vector(to_unsigned(67, 8)),
			5025 => std_logic_vector(to_unsigned(226, 8)),
			5026 => std_logic_vector(to_unsigned(244, 8)),
			5027 => std_logic_vector(to_unsigned(214, 8)),
			5028 => std_logic_vector(to_unsigned(161, 8)),
			5029 => std_logic_vector(to_unsigned(236, 8)),
			5030 => std_logic_vector(to_unsigned(254, 8)),
			5031 => std_logic_vector(to_unsigned(217, 8)),
			5032 => std_logic_vector(to_unsigned(92, 8)),
			5033 => std_logic_vector(to_unsigned(71, 8)),
			5034 => std_logic_vector(to_unsigned(8, 8)),
			5035 => std_logic_vector(to_unsigned(168, 8)),
			5036 => std_logic_vector(to_unsigned(250, 8)),
			5037 => std_logic_vector(to_unsigned(66, 8)),
			5038 => std_logic_vector(to_unsigned(184, 8)),
			5039 => std_logic_vector(to_unsigned(146, 8)),
			5040 => std_logic_vector(to_unsigned(0, 8)),
			5041 => std_logic_vector(to_unsigned(236, 8)),
			5042 => std_logic_vector(to_unsigned(16, 8)),
			5043 => std_logic_vector(to_unsigned(95, 8)),
			5044 => std_logic_vector(to_unsigned(127, 8)),
			5045 => std_logic_vector(to_unsigned(251, 8)),
			5046 => std_logic_vector(to_unsigned(75, 8)),
			5047 => std_logic_vector(to_unsigned(102, 8)),
			5048 => std_logic_vector(to_unsigned(153, 8)),
			5049 => std_logic_vector(to_unsigned(83, 8)),
			5050 => std_logic_vector(to_unsigned(54, 8)),
			5051 => std_logic_vector(to_unsigned(79, 8)),
			5052 => std_logic_vector(to_unsigned(57, 8)),
			5053 => std_logic_vector(to_unsigned(44, 8)),
			5054 => std_logic_vector(to_unsigned(246, 8)),
			5055 => std_logic_vector(to_unsigned(8, 8)),
			5056 => std_logic_vector(to_unsigned(153, 8)),
			5057 => std_logic_vector(to_unsigned(199, 8)),
			5058 => std_logic_vector(to_unsigned(69, 8)),
			5059 => std_logic_vector(to_unsigned(114, 8)),
			5060 => std_logic_vector(to_unsigned(229, 8)),
			5061 => std_logic_vector(to_unsigned(234, 8)),
			5062 => std_logic_vector(to_unsigned(167, 8)),
			5063 => std_logic_vector(to_unsigned(238, 8)),
			5064 => std_logic_vector(to_unsigned(5, 8)),
			5065 => std_logic_vector(to_unsigned(39, 8)),
			5066 => std_logic_vector(to_unsigned(36, 8)),
			5067 => std_logic_vector(to_unsigned(67, 8)),
			5068 => std_logic_vector(to_unsigned(243, 8)),
			5069 => std_logic_vector(to_unsigned(0, 8)),
			5070 => std_logic_vector(to_unsigned(120, 8)),
			5071 => std_logic_vector(to_unsigned(136, 8)),
			5072 => std_logic_vector(to_unsigned(192, 8)),
			5073 => std_logic_vector(to_unsigned(118, 8)),
			5074 => std_logic_vector(to_unsigned(76, 8)),
			5075 => std_logic_vector(to_unsigned(174, 8)),
			5076 => std_logic_vector(to_unsigned(210, 8)),
			5077 => std_logic_vector(to_unsigned(79, 8)),
			5078 => std_logic_vector(to_unsigned(20, 8)),
			5079 => std_logic_vector(to_unsigned(224, 8)),
			5080 => std_logic_vector(to_unsigned(205, 8)),
			5081 => std_logic_vector(to_unsigned(116, 8)),
			5082 => std_logic_vector(to_unsigned(73, 8)),
			5083 => std_logic_vector(to_unsigned(27, 8)),
			5084 => std_logic_vector(to_unsigned(106, 8)),
			5085 => std_logic_vector(to_unsigned(152, 8)),
			5086 => std_logic_vector(to_unsigned(63, 8)),
			5087 => std_logic_vector(to_unsigned(243, 8)),
			5088 => std_logic_vector(to_unsigned(127, 8)),
			5089 => std_logic_vector(to_unsigned(211, 8)),
			5090 => std_logic_vector(to_unsigned(207, 8)),
			5091 => std_logic_vector(to_unsigned(64, 8)),
			5092 => std_logic_vector(to_unsigned(178, 8)),
			5093 => std_logic_vector(to_unsigned(124, 8)),
			5094 => std_logic_vector(to_unsigned(171, 8)),
			5095 => std_logic_vector(to_unsigned(174, 8)),
			5096 => std_logic_vector(to_unsigned(207, 8)),
			5097 => std_logic_vector(to_unsigned(43, 8)),
			5098 => std_logic_vector(to_unsigned(60, 8)),
			5099 => std_logic_vector(to_unsigned(46, 8)),
			5100 => std_logic_vector(to_unsigned(16, 8)),
			5101 => std_logic_vector(to_unsigned(203, 8)),
			5102 => std_logic_vector(to_unsigned(159, 8)),
			5103 => std_logic_vector(to_unsigned(239, 8)),
			5104 => std_logic_vector(to_unsigned(3, 8)),
			5105 => std_logic_vector(to_unsigned(240, 8)),
			5106 => std_logic_vector(to_unsigned(233, 8)),
			5107 => std_logic_vector(to_unsigned(127, 8)),
			5108 => std_logic_vector(to_unsigned(245, 8)),
			5109 => std_logic_vector(to_unsigned(243, 8)),
			5110 => std_logic_vector(to_unsigned(222, 8)),
			5111 => std_logic_vector(to_unsigned(248, 8)),
			5112 => std_logic_vector(to_unsigned(44, 8)),
			5113 => std_logic_vector(to_unsigned(23, 8)),
			5114 => std_logic_vector(to_unsigned(33, 8)),
			5115 => std_logic_vector(to_unsigned(223, 8)),
			5116 => std_logic_vector(to_unsigned(146, 8)),
			5117 => std_logic_vector(to_unsigned(9, 8)),
			5118 => std_logic_vector(to_unsigned(23, 8)),
			5119 => std_logic_vector(to_unsigned(168, 8)),
			5120 => std_logic_vector(to_unsigned(113, 8)),
			5121 => std_logic_vector(to_unsigned(104, 8)),
			5122 => std_logic_vector(to_unsigned(32, 8)),
			5123 => std_logic_vector(to_unsigned(188, 8)),
			5124 => std_logic_vector(to_unsigned(117, 8)),
			5125 => std_logic_vector(to_unsigned(161, 8)),
			5126 => std_logic_vector(to_unsigned(206, 8)),
			5127 => std_logic_vector(to_unsigned(37, 8)),
			5128 => std_logic_vector(to_unsigned(193, 8)),
			5129 => std_logic_vector(to_unsigned(48, 8)),
			5130 => std_logic_vector(to_unsigned(147, 8)),
			5131 => std_logic_vector(to_unsigned(191, 8)),
			5132 => std_logic_vector(to_unsigned(157, 8)),
			5133 => std_logic_vector(to_unsigned(65, 8)),
			5134 => std_logic_vector(to_unsigned(144, 8)),
			5135 => std_logic_vector(to_unsigned(142, 8)),
			5136 => std_logic_vector(to_unsigned(117, 8)),
			5137 => std_logic_vector(to_unsigned(250, 8)),
			5138 => std_logic_vector(to_unsigned(164, 8)),
			5139 => std_logic_vector(to_unsigned(208, 8)),
			5140 => std_logic_vector(to_unsigned(165, 8)),
			5141 => std_logic_vector(to_unsigned(144, 8)),
			5142 => std_logic_vector(to_unsigned(101, 8)),
			5143 => std_logic_vector(to_unsigned(41, 8)),
			5144 => std_logic_vector(to_unsigned(56, 8)),
			5145 => std_logic_vector(to_unsigned(172, 8)),
			5146 => std_logic_vector(to_unsigned(215, 8)),
			5147 => std_logic_vector(to_unsigned(213, 8)),
			5148 => std_logic_vector(to_unsigned(166, 8)),
			5149 => std_logic_vector(to_unsigned(11, 8)),
			5150 => std_logic_vector(to_unsigned(2, 8)),
			5151 => std_logic_vector(to_unsigned(95, 8)),
			5152 => std_logic_vector(to_unsigned(167, 8)),
			5153 => std_logic_vector(to_unsigned(192, 8)),
			5154 => std_logic_vector(to_unsigned(137, 8)),
			5155 => std_logic_vector(to_unsigned(24, 8)),
			5156 => std_logic_vector(to_unsigned(250, 8)),
			5157 => std_logic_vector(to_unsigned(76, 8)),
			5158 => std_logic_vector(to_unsigned(72, 8)),
			5159 => std_logic_vector(to_unsigned(35, 8)),
			5160 => std_logic_vector(to_unsigned(169, 8)),
			5161 => std_logic_vector(to_unsigned(226, 8)),
			5162 => std_logic_vector(to_unsigned(68, 8)),
			5163 => std_logic_vector(to_unsigned(168, 8)),
			5164 => std_logic_vector(to_unsigned(251, 8)),
			5165 => std_logic_vector(to_unsigned(239, 8)),
			5166 => std_logic_vector(to_unsigned(115, 8)),
			5167 => std_logic_vector(to_unsigned(168, 8)),
			5168 => std_logic_vector(to_unsigned(242, 8)),
			5169 => std_logic_vector(to_unsigned(33, 8)),
			5170 => std_logic_vector(to_unsigned(5, 8)),
			5171 => std_logic_vector(to_unsigned(81, 8)),
			5172 => std_logic_vector(to_unsigned(217, 8)),
			5173 => std_logic_vector(to_unsigned(148, 8)),
			5174 => std_logic_vector(to_unsigned(177, 8)),
			5175 => std_logic_vector(to_unsigned(11, 8)),
			5176 => std_logic_vector(to_unsigned(136, 8)),
			5177 => std_logic_vector(to_unsigned(8, 8)),
			5178 => std_logic_vector(to_unsigned(222, 8)),
			5179 => std_logic_vector(to_unsigned(252, 8)),
			5180 => std_logic_vector(to_unsigned(119, 8)),
			5181 => std_logic_vector(to_unsigned(173, 8)),
			5182 => std_logic_vector(to_unsigned(41, 8)),
			5183 => std_logic_vector(to_unsigned(69, 8)),
			5184 => std_logic_vector(to_unsigned(102, 8)),
			5185 => std_logic_vector(to_unsigned(217, 8)),
			5186 => std_logic_vector(to_unsigned(93, 8)),
			5187 => std_logic_vector(to_unsigned(139, 8)),
			5188 => std_logic_vector(to_unsigned(4, 8)),
			5189 => std_logic_vector(to_unsigned(204, 8)),
			5190 => std_logic_vector(to_unsigned(197, 8)),
			5191 => std_logic_vector(to_unsigned(141, 8)),
			5192 => std_logic_vector(to_unsigned(183, 8)),
			5193 => std_logic_vector(to_unsigned(142, 8)),
			5194 => std_logic_vector(to_unsigned(45, 8)),
			5195 => std_logic_vector(to_unsigned(94, 8)),
			5196 => std_logic_vector(to_unsigned(215, 8)),
			5197 => std_logic_vector(to_unsigned(113, 8)),
			5198 => std_logic_vector(to_unsigned(171, 8)),
			5199 => std_logic_vector(to_unsigned(254, 8)),
			5200 => std_logic_vector(to_unsigned(119, 8)),
			5201 => std_logic_vector(to_unsigned(196, 8)),
			5202 => std_logic_vector(to_unsigned(76, 8)),
			5203 => std_logic_vector(to_unsigned(171, 8)),
			5204 => std_logic_vector(to_unsigned(111, 8)),
			5205 => std_logic_vector(to_unsigned(68, 8)),
			5206 => std_logic_vector(to_unsigned(40, 8)),
			5207 => std_logic_vector(to_unsigned(253, 8)),
			5208 => std_logic_vector(to_unsigned(104, 8)),
			5209 => std_logic_vector(to_unsigned(254, 8)),
			5210 => std_logic_vector(to_unsigned(52, 8)),
			5211 => std_logic_vector(to_unsigned(227, 8)),
			5212 => std_logic_vector(to_unsigned(165, 8)),
			5213 => std_logic_vector(to_unsigned(28, 8)),
			5214 => std_logic_vector(to_unsigned(67, 8)),
			5215 => std_logic_vector(to_unsigned(91, 8)),
			5216 => std_logic_vector(to_unsigned(3, 8)),
			5217 => std_logic_vector(to_unsigned(151, 8)),
			5218 => std_logic_vector(to_unsigned(99, 8)),
			5219 => std_logic_vector(to_unsigned(228, 8)),
			5220 => std_logic_vector(to_unsigned(255, 8)),
			5221 => std_logic_vector(to_unsigned(236, 8)),
			5222 => std_logic_vector(to_unsigned(173, 8)),
			5223 => std_logic_vector(to_unsigned(164, 8)),
			5224 => std_logic_vector(to_unsigned(178, 8)),
			5225 => std_logic_vector(to_unsigned(41, 8)),
			5226 => std_logic_vector(to_unsigned(13, 8)),
			5227 => std_logic_vector(to_unsigned(5, 8)),
			5228 => std_logic_vector(to_unsigned(231, 8)),
			5229 => std_logic_vector(to_unsigned(39, 8)),
			5230 => std_logic_vector(to_unsigned(23, 8)),
			5231 => std_logic_vector(to_unsigned(227, 8)),
			5232 => std_logic_vector(to_unsigned(70, 8)),
			5233 => std_logic_vector(to_unsigned(245, 8)),
			5234 => std_logic_vector(to_unsigned(188, 8)),
			5235 => std_logic_vector(to_unsigned(79, 8)),
			5236 => std_logic_vector(to_unsigned(80, 8)),
			5237 => std_logic_vector(to_unsigned(2, 8)),
			5238 => std_logic_vector(to_unsigned(192, 8)),
			5239 => std_logic_vector(to_unsigned(34, 8)),
			5240 => std_logic_vector(to_unsigned(148, 8)),
			5241 => std_logic_vector(to_unsigned(242, 8)),
			5242 => std_logic_vector(to_unsigned(45, 8)),
			5243 => std_logic_vector(to_unsigned(152, 8)),
			5244 => std_logic_vector(to_unsigned(72, 8)),
			5245 => std_logic_vector(to_unsigned(242, 8)),
			5246 => std_logic_vector(to_unsigned(53, 8)),
			5247 => std_logic_vector(to_unsigned(173, 8)),
			5248 => std_logic_vector(to_unsigned(247, 8)),
			5249 => std_logic_vector(to_unsigned(148, 8)),
			5250 => std_logic_vector(to_unsigned(185, 8)),
			5251 => std_logic_vector(to_unsigned(115, 8)),
			5252 => std_logic_vector(to_unsigned(194, 8)),
			5253 => std_logic_vector(to_unsigned(124, 8)),
			5254 => std_logic_vector(to_unsigned(159, 8)),
			5255 => std_logic_vector(to_unsigned(39, 8)),
			5256 => std_logic_vector(to_unsigned(93, 8)),
			5257 => std_logic_vector(to_unsigned(158, 8)),
			5258 => std_logic_vector(to_unsigned(152, 8)),
			5259 => std_logic_vector(to_unsigned(39, 8)),
			5260 => std_logic_vector(to_unsigned(207, 8)),
			5261 => std_logic_vector(to_unsigned(169, 8)),
			5262 => std_logic_vector(to_unsigned(232, 8)),
			5263 => std_logic_vector(to_unsigned(183, 8)),
			5264 => std_logic_vector(to_unsigned(252, 8)),
			5265 => std_logic_vector(to_unsigned(192, 8)),
			5266 => std_logic_vector(to_unsigned(234, 8)),
			5267 => std_logic_vector(to_unsigned(47, 8)),
			5268 => std_logic_vector(to_unsigned(199, 8)),
			5269 => std_logic_vector(to_unsigned(180, 8)),
			5270 => std_logic_vector(to_unsigned(149, 8)),
			5271 => std_logic_vector(to_unsigned(232, 8)),
			5272 => std_logic_vector(to_unsigned(59, 8)),
			5273 => std_logic_vector(to_unsigned(77, 8)),
			5274 => std_logic_vector(to_unsigned(119, 8)),
			5275 => std_logic_vector(to_unsigned(164, 8)),
			5276 => std_logic_vector(to_unsigned(22, 8)),
			5277 => std_logic_vector(to_unsigned(250, 8)),
			5278 => std_logic_vector(to_unsigned(168, 8)),
			5279 => std_logic_vector(to_unsigned(157, 8)),
			5280 => std_logic_vector(to_unsigned(206, 8)),
			5281 => std_logic_vector(to_unsigned(172, 8)),
			5282 => std_logic_vector(to_unsigned(71, 8)),
			5283 => std_logic_vector(to_unsigned(19, 8)),
			5284 => std_logic_vector(to_unsigned(32, 8)),
			5285 => std_logic_vector(to_unsigned(8, 8)),
			5286 => std_logic_vector(to_unsigned(58, 8)),
			5287 => std_logic_vector(to_unsigned(88, 8)),
			5288 => std_logic_vector(to_unsigned(6, 8)),
			5289 => std_logic_vector(to_unsigned(5, 8)),
			5290 => std_logic_vector(to_unsigned(180, 8)),
			5291 => std_logic_vector(to_unsigned(245, 8)),
			5292 => std_logic_vector(to_unsigned(76, 8)),
			5293 => std_logic_vector(to_unsigned(166, 8)),
			5294 => std_logic_vector(to_unsigned(13, 8)),
			5295 => std_logic_vector(to_unsigned(37, 8)),
			5296 => std_logic_vector(to_unsigned(140, 8)),
			5297 => std_logic_vector(to_unsigned(253, 8)),
			5298 => std_logic_vector(to_unsigned(191, 8)),
			5299 => std_logic_vector(to_unsigned(42, 8)),
			5300 => std_logic_vector(to_unsigned(128, 8)),
			5301 => std_logic_vector(to_unsigned(215, 8)),
			5302 => std_logic_vector(to_unsigned(18, 8)),
			5303 => std_logic_vector(to_unsigned(109, 8)),
			5304 => std_logic_vector(to_unsigned(70, 8)),
			5305 => std_logic_vector(to_unsigned(8, 8)),
			5306 => std_logic_vector(to_unsigned(25, 8)),
			5307 => std_logic_vector(to_unsigned(111, 8)),
			5308 => std_logic_vector(to_unsigned(171, 8)),
			5309 => std_logic_vector(to_unsigned(147, 8)),
			5310 => std_logic_vector(to_unsigned(253, 8)),
			5311 => std_logic_vector(to_unsigned(65, 8)),
			5312 => std_logic_vector(to_unsigned(66, 8)),
			5313 => std_logic_vector(to_unsigned(93, 8)),
			5314 => std_logic_vector(to_unsigned(204, 8)),
			5315 => std_logic_vector(to_unsigned(139, 8)),
			5316 => std_logic_vector(to_unsigned(191, 8)),
			5317 => std_logic_vector(to_unsigned(195, 8)),
			5318 => std_logic_vector(to_unsigned(115, 8)),
			5319 => std_logic_vector(to_unsigned(252, 8)),
			5320 => std_logic_vector(to_unsigned(210, 8)),
			5321 => std_logic_vector(to_unsigned(254, 8)),
			5322 => std_logic_vector(to_unsigned(41, 8)),
			5323 => std_logic_vector(to_unsigned(74, 8)),
			5324 => std_logic_vector(to_unsigned(239, 8)),
			5325 => std_logic_vector(to_unsigned(251, 8)),
			5326 => std_logic_vector(to_unsigned(23, 8)),
			5327 => std_logic_vector(to_unsigned(206, 8)),
			5328 => std_logic_vector(to_unsigned(186, 8)),
			5329 => std_logic_vector(to_unsigned(51, 8)),
			5330 => std_logic_vector(to_unsigned(92, 8)),
			5331 => std_logic_vector(to_unsigned(96, 8)),
			5332 => std_logic_vector(to_unsigned(65, 8)),
			5333 => std_logic_vector(to_unsigned(83, 8)),
			5334 => std_logic_vector(to_unsigned(37, 8)),
			5335 => std_logic_vector(to_unsigned(244, 8)),
			5336 => std_logic_vector(to_unsigned(66, 8)),
			5337 => std_logic_vector(to_unsigned(3, 8)),
			5338 => std_logic_vector(to_unsigned(98, 8)),
			5339 => std_logic_vector(to_unsigned(35, 8)),
			5340 => std_logic_vector(to_unsigned(228, 8)),
			5341 => std_logic_vector(to_unsigned(179, 8)),
			5342 => std_logic_vector(to_unsigned(240, 8)),
			5343 => std_logic_vector(to_unsigned(99, 8)),
			5344 => std_logic_vector(to_unsigned(248, 8)),
			5345 => std_logic_vector(to_unsigned(247, 8)),
			5346 => std_logic_vector(to_unsigned(31, 8)),
			5347 => std_logic_vector(to_unsigned(213, 8)),
			5348 => std_logic_vector(to_unsigned(169, 8)),
			5349 => std_logic_vector(to_unsigned(190, 8)),
			5350 => std_logic_vector(to_unsigned(6, 8)),
			5351 => std_logic_vector(to_unsigned(86, 8)),
			5352 => std_logic_vector(to_unsigned(230, 8)),
			5353 => std_logic_vector(to_unsigned(64, 8)),
			5354 => std_logic_vector(to_unsigned(105, 8)),
			5355 => std_logic_vector(to_unsigned(197, 8)),
			5356 => std_logic_vector(to_unsigned(99, 8)),
			5357 => std_logic_vector(to_unsigned(93, 8)),
			5358 => std_logic_vector(to_unsigned(114, 8)),
			5359 => std_logic_vector(to_unsigned(206, 8)),
			5360 => std_logic_vector(to_unsigned(231, 8)),
			5361 => std_logic_vector(to_unsigned(138, 8)),
			5362 => std_logic_vector(to_unsigned(1, 8)),
			5363 => std_logic_vector(to_unsigned(62, 8)),
			5364 => std_logic_vector(to_unsigned(49, 8)),
			5365 => std_logic_vector(to_unsigned(120, 8)),
			5366 => std_logic_vector(to_unsigned(103, 8)),
			5367 => std_logic_vector(to_unsigned(248, 8)),
			5368 => std_logic_vector(to_unsigned(13, 8)),
			5369 => std_logic_vector(to_unsigned(239, 8)),
			5370 => std_logic_vector(to_unsigned(57, 8)),
			5371 => std_logic_vector(to_unsigned(131, 8)),
			5372 => std_logic_vector(to_unsigned(223, 8)),
			5373 => std_logic_vector(to_unsigned(255, 8)),
			5374 => std_logic_vector(to_unsigned(219, 8)),
			5375 => std_logic_vector(to_unsigned(128, 8)),
			5376 => std_logic_vector(to_unsigned(178, 8)),
			5377 => std_logic_vector(to_unsigned(232, 8)),
			5378 => std_logic_vector(to_unsigned(196, 8)),
			5379 => std_logic_vector(to_unsigned(118, 8)),
			5380 => std_logic_vector(to_unsigned(56, 8)),
			5381 => std_logic_vector(to_unsigned(59, 8)),
			5382 => std_logic_vector(to_unsigned(34, 8)),
			5383 => std_logic_vector(to_unsigned(7, 8)),
			5384 => std_logic_vector(to_unsigned(47, 8)),
			5385 => std_logic_vector(to_unsigned(51, 8)),
			5386 => std_logic_vector(to_unsigned(235, 8)),
			5387 => std_logic_vector(to_unsigned(140, 8)),
			5388 => std_logic_vector(to_unsigned(107, 8)),
			5389 => std_logic_vector(to_unsigned(232, 8)),
			5390 => std_logic_vector(to_unsigned(5, 8)),
			5391 => std_logic_vector(to_unsigned(122, 8)),
			5392 => std_logic_vector(to_unsigned(154, 8)),
			5393 => std_logic_vector(to_unsigned(161, 8)),
			5394 => std_logic_vector(to_unsigned(89, 8)),
			5395 => std_logic_vector(to_unsigned(84, 8)),
			5396 => std_logic_vector(to_unsigned(138, 8)),
			5397 => std_logic_vector(to_unsigned(86, 8)),
			5398 => std_logic_vector(to_unsigned(213, 8)),
			5399 => std_logic_vector(to_unsigned(114, 8)),
			5400 => std_logic_vector(to_unsigned(8, 8)),
			5401 => std_logic_vector(to_unsigned(2, 8)),
			5402 => std_logic_vector(to_unsigned(5, 8)),
			5403 => std_logic_vector(to_unsigned(199, 8)),
			5404 => std_logic_vector(to_unsigned(101, 8)),
			5405 => std_logic_vector(to_unsigned(113, 8)),
			5406 => std_logic_vector(to_unsigned(126, 8)),
			5407 => std_logic_vector(to_unsigned(27, 8)),
			5408 => std_logic_vector(to_unsigned(131, 8)),
			5409 => std_logic_vector(to_unsigned(130, 8)),
			5410 => std_logic_vector(to_unsigned(169, 8)),
			5411 => std_logic_vector(to_unsigned(183, 8)),
			5412 => std_logic_vector(to_unsigned(130, 8)),
			5413 => std_logic_vector(to_unsigned(73, 8)),
			5414 => std_logic_vector(to_unsigned(175, 8)),
			5415 => std_logic_vector(to_unsigned(49, 8)),
			5416 => std_logic_vector(to_unsigned(92, 8)),
			5417 => std_logic_vector(to_unsigned(150, 8)),
			5418 => std_logic_vector(to_unsigned(209, 8)),
			5419 => std_logic_vector(to_unsigned(23, 8)),
			5420 => std_logic_vector(to_unsigned(135, 8)),
			5421 => std_logic_vector(to_unsigned(190, 8)),
			5422 => std_logic_vector(to_unsigned(67, 8)),
			5423 => std_logic_vector(to_unsigned(68, 8)),
			5424 => std_logic_vector(to_unsigned(69, 8)),
			5425 => std_logic_vector(to_unsigned(153, 8)),
			5426 => std_logic_vector(to_unsigned(26, 8)),
			5427 => std_logic_vector(to_unsigned(96, 8)),
			5428 => std_logic_vector(to_unsigned(182, 8)),
			5429 => std_logic_vector(to_unsigned(171, 8)),
			5430 => std_logic_vector(to_unsigned(80, 8)),
			5431 => std_logic_vector(to_unsigned(162, 8)),
			5432 => std_logic_vector(to_unsigned(86, 8)),
			5433 => std_logic_vector(to_unsigned(65, 8)),
			5434 => std_logic_vector(to_unsigned(27, 8)),
			5435 => std_logic_vector(to_unsigned(63, 8)),
			5436 => std_logic_vector(to_unsigned(172, 8)),
			5437 => std_logic_vector(to_unsigned(45, 8)),
			5438 => std_logic_vector(to_unsigned(171, 8)),
			5439 => std_logic_vector(to_unsigned(199, 8)),
			5440 => std_logic_vector(to_unsigned(7, 8)),
			5441 => std_logic_vector(to_unsigned(2, 8)),
			5442 => std_logic_vector(to_unsigned(56, 8)),
			5443 => std_logic_vector(to_unsigned(206, 8)),
			5444 => std_logic_vector(to_unsigned(217, 8)),
			5445 => std_logic_vector(to_unsigned(162, 8)),
			5446 => std_logic_vector(to_unsigned(224, 8)),
			5447 => std_logic_vector(to_unsigned(239, 8)),
			5448 => std_logic_vector(to_unsigned(36, 8)),
			5449 => std_logic_vector(to_unsigned(46, 8)),
			5450 => std_logic_vector(to_unsigned(93, 8)),
			5451 => std_logic_vector(to_unsigned(10, 8)),
			5452 => std_logic_vector(to_unsigned(34, 8)),
			5453 => std_logic_vector(to_unsigned(120, 8)),
			5454 => std_logic_vector(to_unsigned(159, 8)),
			5455 => std_logic_vector(to_unsigned(229, 8)),
			5456 => std_logic_vector(to_unsigned(170, 8)),
			5457 => std_logic_vector(to_unsigned(139, 8)),
			5458 => std_logic_vector(to_unsigned(72, 8)),
			5459 => std_logic_vector(to_unsigned(208, 8)),
			5460 => std_logic_vector(to_unsigned(151, 8)),
			5461 => std_logic_vector(to_unsigned(164, 8)),
			5462 => std_logic_vector(to_unsigned(27, 8)),
			5463 => std_logic_vector(to_unsigned(2, 8)),
			5464 => std_logic_vector(to_unsigned(122, 8)),
			5465 => std_logic_vector(to_unsigned(175, 8)),
			5466 => std_logic_vector(to_unsigned(9, 8)),
			5467 => std_logic_vector(to_unsigned(105, 8)),
			5468 => std_logic_vector(to_unsigned(232, 8)),
			5469 => std_logic_vector(to_unsigned(221, 8)),
			5470 => std_logic_vector(to_unsigned(153, 8)),
			5471 => std_logic_vector(to_unsigned(229, 8)),
			5472 => std_logic_vector(to_unsigned(242, 8)),
			5473 => std_logic_vector(to_unsigned(128, 8)),
			5474 => std_logic_vector(to_unsigned(177, 8)),
			5475 => std_logic_vector(to_unsigned(225, 8)),
			5476 => std_logic_vector(to_unsigned(103, 8)),
			5477 => std_logic_vector(to_unsigned(173, 8)),
			5478 => std_logic_vector(to_unsigned(201, 8)),
			5479 => std_logic_vector(to_unsigned(110, 8)),
			5480 => std_logic_vector(to_unsigned(156, 8)),
			5481 => std_logic_vector(to_unsigned(177, 8)),
			5482 => std_logic_vector(to_unsigned(133, 8)),
			5483 => std_logic_vector(to_unsigned(88, 8)),
			5484 => std_logic_vector(to_unsigned(45, 8)),
			5485 => std_logic_vector(to_unsigned(16, 8)),
			5486 => std_logic_vector(to_unsigned(254, 8)),
			5487 => std_logic_vector(to_unsigned(29, 8)),
			5488 => std_logic_vector(to_unsigned(16, 8)),
			5489 => std_logic_vector(to_unsigned(10, 8)),
			5490 => std_logic_vector(to_unsigned(43, 8)),
			5491 => std_logic_vector(to_unsigned(211, 8)),
			5492 => std_logic_vector(to_unsigned(105, 8)),
			5493 => std_logic_vector(to_unsigned(223, 8)),
			5494 => std_logic_vector(to_unsigned(205, 8)),
			5495 => std_logic_vector(to_unsigned(9, 8)),
			5496 => std_logic_vector(to_unsigned(169, 8)),
			5497 => std_logic_vector(to_unsigned(7, 8)),
			5498 => std_logic_vector(to_unsigned(224, 8)),
			5499 => std_logic_vector(to_unsigned(19, 8)),
			5500 => std_logic_vector(to_unsigned(83, 8)),
			5501 => std_logic_vector(to_unsigned(28, 8)),
			5502 => std_logic_vector(to_unsigned(116, 8)),
			5503 => std_logic_vector(to_unsigned(155, 8)),
			5504 => std_logic_vector(to_unsigned(58, 8)),
			5505 => std_logic_vector(to_unsigned(122, 8)),
			5506 => std_logic_vector(to_unsigned(214, 8)),
			5507 => std_logic_vector(to_unsigned(47, 8)),
			5508 => std_logic_vector(to_unsigned(48, 8)),
			5509 => std_logic_vector(to_unsigned(68, 8)),
			5510 => std_logic_vector(to_unsigned(145, 8)),
			5511 => std_logic_vector(to_unsigned(15, 8)),
			5512 => std_logic_vector(to_unsigned(215, 8)),
			5513 => std_logic_vector(to_unsigned(93, 8)),
			5514 => std_logic_vector(to_unsigned(92, 8)),
			5515 => std_logic_vector(to_unsigned(93, 8)),
			5516 => std_logic_vector(to_unsigned(26, 8)),
			5517 => std_logic_vector(to_unsigned(199, 8)),
			5518 => std_logic_vector(to_unsigned(141, 8)),
			5519 => std_logic_vector(to_unsigned(14, 8)),
			5520 => std_logic_vector(to_unsigned(79, 8)),
			5521 => std_logic_vector(to_unsigned(6, 8)),
			5522 => std_logic_vector(to_unsigned(2, 8)),
			5523 => std_logic_vector(to_unsigned(175, 8)),
			5524 => std_logic_vector(to_unsigned(52, 8)),
			5525 => std_logic_vector(to_unsigned(30, 8)),
			5526 => std_logic_vector(to_unsigned(72, 8)),
			5527 => std_logic_vector(to_unsigned(94, 8)),
			5528 => std_logic_vector(to_unsigned(77, 8)),
			5529 => std_logic_vector(to_unsigned(210, 8)),
			5530 => std_logic_vector(to_unsigned(154, 8)),
			5531 => std_logic_vector(to_unsigned(17, 8)),
			5532 => std_logic_vector(to_unsigned(207, 8)),
			5533 => std_logic_vector(to_unsigned(107, 8)),
			5534 => std_logic_vector(to_unsigned(131, 8)),
			5535 => std_logic_vector(to_unsigned(163, 8)),
			5536 => std_logic_vector(to_unsigned(254, 8)),
			5537 => std_logic_vector(to_unsigned(120, 8)),
			5538 => std_logic_vector(to_unsigned(48, 8)),
			5539 => std_logic_vector(to_unsigned(130, 8)),
			5540 => std_logic_vector(to_unsigned(156, 8)),
			5541 => std_logic_vector(to_unsigned(226, 8)),
			5542 => std_logic_vector(to_unsigned(184, 8)),
			5543 => std_logic_vector(to_unsigned(37, 8)),
			5544 => std_logic_vector(to_unsigned(170, 8)),
			5545 => std_logic_vector(to_unsigned(131, 8)),
			5546 => std_logic_vector(to_unsigned(125, 8)),
			5547 => std_logic_vector(to_unsigned(82, 8)),
			5548 => std_logic_vector(to_unsigned(78, 8)),
			5549 => std_logic_vector(to_unsigned(23, 8)),
			5550 => std_logic_vector(to_unsigned(154, 8)),
			5551 => std_logic_vector(to_unsigned(11, 8)),
			5552 => std_logic_vector(to_unsigned(238, 8)),
			5553 => std_logic_vector(to_unsigned(95, 8)),
			5554 => std_logic_vector(to_unsigned(25, 8)),
			5555 => std_logic_vector(to_unsigned(249, 8)),
			5556 => std_logic_vector(to_unsigned(225, 8)),
			5557 => std_logic_vector(to_unsigned(4, 8)),
			5558 => std_logic_vector(to_unsigned(237, 8)),
			5559 => std_logic_vector(to_unsigned(89, 8)),
			5560 => std_logic_vector(to_unsigned(80, 8)),
			5561 => std_logic_vector(to_unsigned(202, 8)),
			5562 => std_logic_vector(to_unsigned(134, 8)),
			5563 => std_logic_vector(to_unsigned(12, 8)),
			5564 => std_logic_vector(to_unsigned(194, 8)),
			5565 => std_logic_vector(to_unsigned(35, 8)),
			5566 => std_logic_vector(to_unsigned(96, 8)),
			5567 => std_logic_vector(to_unsigned(44, 8)),
			5568 => std_logic_vector(to_unsigned(197, 8)),
			5569 => std_logic_vector(to_unsigned(110, 8)),
			5570 => std_logic_vector(to_unsigned(129, 8)),
			5571 => std_logic_vector(to_unsigned(251, 8)),
			5572 => std_logic_vector(to_unsigned(197, 8)),
			5573 => std_logic_vector(to_unsigned(9, 8)),
			5574 => std_logic_vector(to_unsigned(44, 8)),
			5575 => std_logic_vector(to_unsigned(209, 8)),
			5576 => std_logic_vector(to_unsigned(192, 8)),
			5577 => std_logic_vector(to_unsigned(223, 8)),
			5578 => std_logic_vector(to_unsigned(124, 8)),
			5579 => std_logic_vector(to_unsigned(130, 8)),
			5580 => std_logic_vector(to_unsigned(240, 8)),
			5581 => std_logic_vector(to_unsigned(247, 8)),
			5582 => std_logic_vector(to_unsigned(119, 8)),
			5583 => std_logic_vector(to_unsigned(9, 8)),
			5584 => std_logic_vector(to_unsigned(233, 8)),
			5585 => std_logic_vector(to_unsigned(19, 8)),
			5586 => std_logic_vector(to_unsigned(210, 8)),
			5587 => std_logic_vector(to_unsigned(79, 8)),
			5588 => std_logic_vector(to_unsigned(110, 8)),
			5589 => std_logic_vector(to_unsigned(234, 8)),
			5590 => std_logic_vector(to_unsigned(120, 8)),
			5591 => std_logic_vector(to_unsigned(224, 8)),
			5592 => std_logic_vector(to_unsigned(130, 8)),
			5593 => std_logic_vector(to_unsigned(193, 8)),
			5594 => std_logic_vector(to_unsigned(129, 8)),
			5595 => std_logic_vector(to_unsigned(0, 8)),
			5596 => std_logic_vector(to_unsigned(37, 8)),
			5597 => std_logic_vector(to_unsigned(5, 8)),
			5598 => std_logic_vector(to_unsigned(133, 8)),
			5599 => std_logic_vector(to_unsigned(225, 8)),
			5600 => std_logic_vector(to_unsigned(136, 8)),
			5601 => std_logic_vector(to_unsigned(52, 8)),
			5602 => std_logic_vector(to_unsigned(141, 8)),
			5603 => std_logic_vector(to_unsigned(152, 8)),
			5604 => std_logic_vector(to_unsigned(233, 8)),
			5605 => std_logic_vector(to_unsigned(145, 8)),
			5606 => std_logic_vector(to_unsigned(222, 8)),
			5607 => std_logic_vector(to_unsigned(127, 8)),
			5608 => std_logic_vector(to_unsigned(193, 8)),
			5609 => std_logic_vector(to_unsigned(101, 8)),
			5610 => std_logic_vector(to_unsigned(127, 8)),
			5611 => std_logic_vector(to_unsigned(84, 8)),
			5612 => std_logic_vector(to_unsigned(161, 8)),
			5613 => std_logic_vector(to_unsigned(12, 8)),
			5614 => std_logic_vector(to_unsigned(242, 8)),
			5615 => std_logic_vector(to_unsigned(72, 8)),
			5616 => std_logic_vector(to_unsigned(148, 8)),
			5617 => std_logic_vector(to_unsigned(137, 8)),
			5618 => std_logic_vector(to_unsigned(186, 8)),
			5619 => std_logic_vector(to_unsigned(55, 8)),
			5620 => std_logic_vector(to_unsigned(176, 8)),
			5621 => std_logic_vector(to_unsigned(162, 8)),
			5622 => std_logic_vector(to_unsigned(128, 8)),
			5623 => std_logic_vector(to_unsigned(203, 8)),
			5624 => std_logic_vector(to_unsigned(84, 8)),
			5625 => std_logic_vector(to_unsigned(229, 8)),
			5626 => std_logic_vector(to_unsigned(21, 8)),
			5627 => std_logic_vector(to_unsigned(223, 8)),
			5628 => std_logic_vector(to_unsigned(61, 8)),
			5629 => std_logic_vector(to_unsigned(74, 8)),
			5630 => std_logic_vector(to_unsigned(84, 8)),
			5631 => std_logic_vector(to_unsigned(46, 8)),
			5632 => std_logic_vector(to_unsigned(93, 8)),
			5633 => std_logic_vector(to_unsigned(14, 8)),
			5634 => std_logic_vector(to_unsigned(219, 8)),
			5635 => std_logic_vector(to_unsigned(201, 8)),
			5636 => std_logic_vector(to_unsigned(246, 8)),
			5637 => std_logic_vector(to_unsigned(191, 8)),
			5638 => std_logic_vector(to_unsigned(190, 8)),
			5639 => std_logic_vector(to_unsigned(53, 8)),
			5640 => std_logic_vector(to_unsigned(195, 8)),
			5641 => std_logic_vector(to_unsigned(21, 8)),
			5642 => std_logic_vector(to_unsigned(213, 8)),
			5643 => std_logic_vector(to_unsigned(160, 8)),
			5644 => std_logic_vector(to_unsigned(176, 8)),
			5645 => std_logic_vector(to_unsigned(10, 8)),
			5646 => std_logic_vector(to_unsigned(176, 8)),
			5647 => std_logic_vector(to_unsigned(109, 8)),
			5648 => std_logic_vector(to_unsigned(74, 8)),
			5649 => std_logic_vector(to_unsigned(11, 8)),
			5650 => std_logic_vector(to_unsigned(219, 8)),
			5651 => std_logic_vector(to_unsigned(7, 8)),
			5652 => std_logic_vector(to_unsigned(146, 8)),
			5653 => std_logic_vector(to_unsigned(245, 8)),
			5654 => std_logic_vector(to_unsigned(59, 8)),
			5655 => std_logic_vector(to_unsigned(13, 8)),
			5656 => std_logic_vector(to_unsigned(55, 8)),
			5657 => std_logic_vector(to_unsigned(40, 8)),
			5658 => std_logic_vector(to_unsigned(245, 8)),
			5659 => std_logic_vector(to_unsigned(105, 8)),
			5660 => std_logic_vector(to_unsigned(198, 8)),
			5661 => std_logic_vector(to_unsigned(197, 8)),
			5662 => std_logic_vector(to_unsigned(247, 8)),
			5663 => std_logic_vector(to_unsigned(72, 8)),
			5664 => std_logic_vector(to_unsigned(141, 8)),
			5665 => std_logic_vector(to_unsigned(191, 8)),
			5666 => std_logic_vector(to_unsigned(151, 8)),
			5667 => std_logic_vector(to_unsigned(87, 8)),
			5668 => std_logic_vector(to_unsigned(10, 8)),
			5669 => std_logic_vector(to_unsigned(153, 8)),
			5670 => std_logic_vector(to_unsigned(39, 8)),
			5671 => std_logic_vector(to_unsigned(237, 8)),
			5672 => std_logic_vector(to_unsigned(25, 8)),
			5673 => std_logic_vector(to_unsigned(33, 8)),
			5674 => std_logic_vector(to_unsigned(94, 8)),
			5675 => std_logic_vector(to_unsigned(245, 8)),
			5676 => std_logic_vector(to_unsigned(148, 8)),
			5677 => std_logic_vector(to_unsigned(215, 8)),
			5678 => std_logic_vector(to_unsigned(4, 8)),
			5679 => std_logic_vector(to_unsigned(97, 8)),
			5680 => std_logic_vector(to_unsigned(112, 8)),
			5681 => std_logic_vector(to_unsigned(222, 8)),
			5682 => std_logic_vector(to_unsigned(57, 8)),
			5683 => std_logic_vector(to_unsigned(232, 8)),
			5684 => std_logic_vector(to_unsigned(168, 8)),
			5685 => std_logic_vector(to_unsigned(244, 8)),
			5686 => std_logic_vector(to_unsigned(199, 8)),
			5687 => std_logic_vector(to_unsigned(214, 8)),
			5688 => std_logic_vector(to_unsigned(224, 8)),
			5689 => std_logic_vector(to_unsigned(230, 8)),
			5690 => std_logic_vector(to_unsigned(24, 8)),
			5691 => std_logic_vector(to_unsigned(94, 8)),
			5692 => std_logic_vector(to_unsigned(170, 8)),
			5693 => std_logic_vector(to_unsigned(203, 8)),
			5694 => std_logic_vector(to_unsigned(113, 8)),
			5695 => std_logic_vector(to_unsigned(146, 8)),
			5696 => std_logic_vector(to_unsigned(109, 8)),
			5697 => std_logic_vector(to_unsigned(1, 8)),
			5698 => std_logic_vector(to_unsigned(60, 8)),
			5699 => std_logic_vector(to_unsigned(29, 8)),
			5700 => std_logic_vector(to_unsigned(201, 8)),
			5701 => std_logic_vector(to_unsigned(45, 8)),
			5702 => std_logic_vector(to_unsigned(92, 8)),
			5703 => std_logic_vector(to_unsigned(92, 8)),
			5704 => std_logic_vector(to_unsigned(250, 8)),
			5705 => std_logic_vector(to_unsigned(118, 8)),
			5706 => std_logic_vector(to_unsigned(94, 8)),
			5707 => std_logic_vector(to_unsigned(12, 8)),
			5708 => std_logic_vector(to_unsigned(244, 8)),
			5709 => std_logic_vector(to_unsigned(254, 8)),
			5710 => std_logic_vector(to_unsigned(137, 8)),
			5711 => std_logic_vector(to_unsigned(50, 8)),
			5712 => std_logic_vector(to_unsigned(54, 8)),
			5713 => std_logic_vector(to_unsigned(235, 8)),
			5714 => std_logic_vector(to_unsigned(71, 8)),
			5715 => std_logic_vector(to_unsigned(137, 8)),
			5716 => std_logic_vector(to_unsigned(247, 8)),
			5717 => std_logic_vector(to_unsigned(196, 8)),
			5718 => std_logic_vector(to_unsigned(234, 8)),
			5719 => std_logic_vector(to_unsigned(162, 8)),
			5720 => std_logic_vector(to_unsigned(42, 8)),
			5721 => std_logic_vector(to_unsigned(133, 8)),
			5722 => std_logic_vector(to_unsigned(188, 8)),
			5723 => std_logic_vector(to_unsigned(195, 8)),
			5724 => std_logic_vector(to_unsigned(220, 8)),
			5725 => std_logic_vector(to_unsigned(171, 8)),
			5726 => std_logic_vector(to_unsigned(88, 8)),
			5727 => std_logic_vector(to_unsigned(181, 8)),
			5728 => std_logic_vector(to_unsigned(176, 8)),
			5729 => std_logic_vector(to_unsigned(228, 8)),
			5730 => std_logic_vector(to_unsigned(57, 8)),
			5731 => std_logic_vector(to_unsigned(96, 8)),
			5732 => std_logic_vector(to_unsigned(8, 8)),
			5733 => std_logic_vector(to_unsigned(0, 8)),
			5734 => std_logic_vector(to_unsigned(156, 8)),
			5735 => std_logic_vector(to_unsigned(125, 8)),
			5736 => std_logic_vector(to_unsigned(2, 8)),
			5737 => std_logic_vector(to_unsigned(75, 8)),
			5738 => std_logic_vector(to_unsigned(157, 8)),
			5739 => std_logic_vector(to_unsigned(58, 8)),
			5740 => std_logic_vector(to_unsigned(90, 8)),
			5741 => std_logic_vector(to_unsigned(37, 8)),
			5742 => std_logic_vector(to_unsigned(142, 8)),
			5743 => std_logic_vector(to_unsigned(194, 8)),
			5744 => std_logic_vector(to_unsigned(40, 8)),
			5745 => std_logic_vector(to_unsigned(96, 8)),
			5746 => std_logic_vector(to_unsigned(121, 8)),
			5747 => std_logic_vector(to_unsigned(57, 8)),
			5748 => std_logic_vector(to_unsigned(240, 8)),
			5749 => std_logic_vector(to_unsigned(226, 8)),
			5750 => std_logic_vector(to_unsigned(84, 8)),
			5751 => std_logic_vector(to_unsigned(208, 8)),
			5752 => std_logic_vector(to_unsigned(169, 8)),
			5753 => std_logic_vector(to_unsigned(74, 8)),
			5754 => std_logic_vector(to_unsigned(239, 8)),
			5755 => std_logic_vector(to_unsigned(212, 8)),
			5756 => std_logic_vector(to_unsigned(161, 8)),
			5757 => std_logic_vector(to_unsigned(43, 8)),
			5758 => std_logic_vector(to_unsigned(54, 8)),
			5759 => std_logic_vector(to_unsigned(176, 8)),
			5760 => std_logic_vector(to_unsigned(66, 8)),
			5761 => std_logic_vector(to_unsigned(107, 8)),
			5762 => std_logic_vector(to_unsigned(85, 8)),
			5763 => std_logic_vector(to_unsigned(117, 8)),
			5764 => std_logic_vector(to_unsigned(243, 8)),
			5765 => std_logic_vector(to_unsigned(245, 8)),
			5766 => std_logic_vector(to_unsigned(168, 8)),
			5767 => std_logic_vector(to_unsigned(150, 8)),
			5768 => std_logic_vector(to_unsigned(130, 8)),
			5769 => std_logic_vector(to_unsigned(19, 8)),
			5770 => std_logic_vector(to_unsigned(220, 8)),
			5771 => std_logic_vector(to_unsigned(121, 8)),
			5772 => std_logic_vector(to_unsigned(24, 8)),
			5773 => std_logic_vector(to_unsigned(13, 8)),
			5774 => std_logic_vector(to_unsigned(163, 8)),
			5775 => std_logic_vector(to_unsigned(235, 8)),
			5776 => std_logic_vector(to_unsigned(44, 8)),
			5777 => std_logic_vector(to_unsigned(168, 8)),
			5778 => std_logic_vector(to_unsigned(66, 8)),
			5779 => std_logic_vector(to_unsigned(63, 8)),
			5780 => std_logic_vector(to_unsigned(187, 8)),
			5781 => std_logic_vector(to_unsigned(26, 8)),
			5782 => std_logic_vector(to_unsigned(212, 8)),
			5783 => std_logic_vector(to_unsigned(58, 8)),
			5784 => std_logic_vector(to_unsigned(2, 8)),
			5785 => std_logic_vector(to_unsigned(6, 8)),
			5786 => std_logic_vector(to_unsigned(185, 8)),
			5787 => std_logic_vector(to_unsigned(183, 8)),
			5788 => std_logic_vector(to_unsigned(253, 8)),
			5789 => std_logic_vector(to_unsigned(93, 8)),
			5790 => std_logic_vector(to_unsigned(189, 8)),
			5791 => std_logic_vector(to_unsigned(187, 8)),
			5792 => std_logic_vector(to_unsigned(222, 8)),
			5793 => std_logic_vector(to_unsigned(73, 8)),
			5794 => std_logic_vector(to_unsigned(130, 8)),
			5795 => std_logic_vector(to_unsigned(234, 8)),
			5796 => std_logic_vector(to_unsigned(203, 8)),
			5797 => std_logic_vector(to_unsigned(25, 8)),
			5798 => std_logic_vector(to_unsigned(215, 8)),
			5799 => std_logic_vector(to_unsigned(43, 8)),
			5800 => std_logic_vector(to_unsigned(7, 8)),
			5801 => std_logic_vector(to_unsigned(115, 8)),
			5802 => std_logic_vector(to_unsigned(196, 8)),
			5803 => std_logic_vector(to_unsigned(68, 8)),
			5804 => std_logic_vector(to_unsigned(9, 8)),
			5805 => std_logic_vector(to_unsigned(162, 8)),
			5806 => std_logic_vector(to_unsigned(129, 8)),
			5807 => std_logic_vector(to_unsigned(165, 8)),
			5808 => std_logic_vector(to_unsigned(48, 8)),
			5809 => std_logic_vector(to_unsigned(140, 8)),
			5810 => std_logic_vector(to_unsigned(11, 8)),
			5811 => std_logic_vector(to_unsigned(184, 8)),
			5812 => std_logic_vector(to_unsigned(100, 8)),
			5813 => std_logic_vector(to_unsigned(201, 8)),
			5814 => std_logic_vector(to_unsigned(61, 8)),
			5815 => std_logic_vector(to_unsigned(240, 8)),
			5816 => std_logic_vector(to_unsigned(71, 8)),
			5817 => std_logic_vector(to_unsigned(15, 8)),
			5818 => std_logic_vector(to_unsigned(72, 8)),
			5819 => std_logic_vector(to_unsigned(120, 8)),
			5820 => std_logic_vector(to_unsigned(184, 8)),
			5821 => std_logic_vector(to_unsigned(173, 8)),
			5822 => std_logic_vector(to_unsigned(21, 8)),
			5823 => std_logic_vector(to_unsigned(109, 8)),
			5824 => std_logic_vector(to_unsigned(64, 8)),
			5825 => std_logic_vector(to_unsigned(92, 8)),
			5826 => std_logic_vector(to_unsigned(32, 8)),
			5827 => std_logic_vector(to_unsigned(237, 8)),
			5828 => std_logic_vector(to_unsigned(87, 8)),
			5829 => std_logic_vector(to_unsigned(234, 8)),
			5830 => std_logic_vector(to_unsigned(176, 8)),
			5831 => std_logic_vector(to_unsigned(208, 8)),
			5832 => std_logic_vector(to_unsigned(13, 8)),
			5833 => std_logic_vector(to_unsigned(46, 8)),
			5834 => std_logic_vector(to_unsigned(247, 8)),
			5835 => std_logic_vector(to_unsigned(80, 8)),
			5836 => std_logic_vector(to_unsigned(212, 8)),
			5837 => std_logic_vector(to_unsigned(29, 8)),
			5838 => std_logic_vector(to_unsigned(182, 8)),
			5839 => std_logic_vector(to_unsigned(38, 8)),
			5840 => std_logic_vector(to_unsigned(227, 8)),
			5841 => std_logic_vector(to_unsigned(66, 8)),
			5842 => std_logic_vector(to_unsigned(72, 8)),
			5843 => std_logic_vector(to_unsigned(215, 8)),
			5844 => std_logic_vector(to_unsigned(3, 8)),
			5845 => std_logic_vector(to_unsigned(87, 8)),
			5846 => std_logic_vector(to_unsigned(22, 8)),
			5847 => std_logic_vector(to_unsigned(132, 8)),
			5848 => std_logic_vector(to_unsigned(118, 8)),
			5849 => std_logic_vector(to_unsigned(104, 8)),
			5850 => std_logic_vector(to_unsigned(141, 8)),
			5851 => std_logic_vector(to_unsigned(42, 8)),
			5852 => std_logic_vector(to_unsigned(138, 8)),
			5853 => std_logic_vector(to_unsigned(214, 8)),
			5854 => std_logic_vector(to_unsigned(9, 8)),
			5855 => std_logic_vector(to_unsigned(67, 8)),
			5856 => std_logic_vector(to_unsigned(172, 8)),
			5857 => std_logic_vector(to_unsigned(25, 8)),
			5858 => std_logic_vector(to_unsigned(46, 8)),
			5859 => std_logic_vector(to_unsigned(244, 8)),
			5860 => std_logic_vector(to_unsigned(222, 8)),
			5861 => std_logic_vector(to_unsigned(51, 8)),
			5862 => std_logic_vector(to_unsigned(167, 8)),
			5863 => std_logic_vector(to_unsigned(54, 8)),
			5864 => std_logic_vector(to_unsigned(54, 8)),
			5865 => std_logic_vector(to_unsigned(167, 8)),
			5866 => std_logic_vector(to_unsigned(136, 8)),
			5867 => std_logic_vector(to_unsigned(73, 8)),
			5868 => std_logic_vector(to_unsigned(250, 8)),
			5869 => std_logic_vector(to_unsigned(40, 8)),
			5870 => std_logic_vector(to_unsigned(127, 8)),
			5871 => std_logic_vector(to_unsigned(53, 8)),
			5872 => std_logic_vector(to_unsigned(166, 8)),
			5873 => std_logic_vector(to_unsigned(225, 8)),
			5874 => std_logic_vector(to_unsigned(18, 8)),
			5875 => std_logic_vector(to_unsigned(185, 8)),
			5876 => std_logic_vector(to_unsigned(42, 8)),
			5877 => std_logic_vector(to_unsigned(44, 8)),
			5878 => std_logic_vector(to_unsigned(175, 8)),
			5879 => std_logic_vector(to_unsigned(96, 8)),
			5880 => std_logic_vector(to_unsigned(8, 8)),
			5881 => std_logic_vector(to_unsigned(93, 8)),
			5882 => std_logic_vector(to_unsigned(31, 8)),
			5883 => std_logic_vector(to_unsigned(128, 8)),
			5884 => std_logic_vector(to_unsigned(93, 8)),
			5885 => std_logic_vector(to_unsigned(175, 8)),
			5886 => std_logic_vector(to_unsigned(167, 8)),
			5887 => std_logic_vector(to_unsigned(238, 8)),
			5888 => std_logic_vector(to_unsigned(48, 8)),
			5889 => std_logic_vector(to_unsigned(61, 8)),
			5890 => std_logic_vector(to_unsigned(87, 8)),
			5891 => std_logic_vector(to_unsigned(173, 8)),
			5892 => std_logic_vector(to_unsigned(219, 8)),
			5893 => std_logic_vector(to_unsigned(119, 8)),
			5894 => std_logic_vector(to_unsigned(37, 8)),
			5895 => std_logic_vector(to_unsigned(176, 8)),
			5896 => std_logic_vector(to_unsigned(112, 8)),
			5897 => std_logic_vector(to_unsigned(122, 8)),
			5898 => std_logic_vector(to_unsigned(15, 8)),
			5899 => std_logic_vector(to_unsigned(155, 8)),
			5900 => std_logic_vector(to_unsigned(243, 8)),
			5901 => std_logic_vector(to_unsigned(211, 8)),
			5902 => std_logic_vector(to_unsigned(242, 8)),
			5903 => std_logic_vector(to_unsigned(107, 8)),
			5904 => std_logic_vector(to_unsigned(141, 8)),
			5905 => std_logic_vector(to_unsigned(236, 8)),
			5906 => std_logic_vector(to_unsigned(154, 8)),
			5907 => std_logic_vector(to_unsigned(242, 8)),
			5908 => std_logic_vector(to_unsigned(77, 8)),
			5909 => std_logic_vector(to_unsigned(224, 8)),
			5910 => std_logic_vector(to_unsigned(46, 8)),
			5911 => std_logic_vector(to_unsigned(42, 8)),
			5912 => std_logic_vector(to_unsigned(219, 8)),
			5913 => std_logic_vector(to_unsigned(140, 8)),
			5914 => std_logic_vector(to_unsigned(105, 8)),
			5915 => std_logic_vector(to_unsigned(113, 8)),
			5916 => std_logic_vector(to_unsigned(159, 8)),
			5917 => std_logic_vector(to_unsigned(76, 8)),
			5918 => std_logic_vector(to_unsigned(58, 8)),
			5919 => std_logic_vector(to_unsigned(222, 8)),
			5920 => std_logic_vector(to_unsigned(107, 8)),
			5921 => std_logic_vector(to_unsigned(132, 8)),
			5922 => std_logic_vector(to_unsigned(80, 8)),
			5923 => std_logic_vector(to_unsigned(122, 8)),
			5924 => std_logic_vector(to_unsigned(75, 8)),
			5925 => std_logic_vector(to_unsigned(103, 8)),
			5926 => std_logic_vector(to_unsigned(74, 8)),
			5927 => std_logic_vector(to_unsigned(110, 8)),
			5928 => std_logic_vector(to_unsigned(145, 8)),
			5929 => std_logic_vector(to_unsigned(27, 8)),
			5930 => std_logic_vector(to_unsigned(224, 8)),
			5931 => std_logic_vector(to_unsigned(95, 8)),
			5932 => std_logic_vector(to_unsigned(227, 8)),
			5933 => std_logic_vector(to_unsigned(216, 8)),
			5934 => std_logic_vector(to_unsigned(99, 8)),
			5935 => std_logic_vector(to_unsigned(181, 8)),
			5936 => std_logic_vector(to_unsigned(148, 8)),
			5937 => std_logic_vector(to_unsigned(149, 8)),
			5938 => std_logic_vector(to_unsigned(122, 8)),
			5939 => std_logic_vector(to_unsigned(78, 8)),
			5940 => std_logic_vector(to_unsigned(42, 8)),
			5941 => std_logic_vector(to_unsigned(146, 8)),
			5942 => std_logic_vector(to_unsigned(191, 8)),
			5943 => std_logic_vector(to_unsigned(183, 8)),
			5944 => std_logic_vector(to_unsigned(104, 8)),
			5945 => std_logic_vector(to_unsigned(248, 8)),
			5946 => std_logic_vector(to_unsigned(140, 8)),
			5947 => std_logic_vector(to_unsigned(162, 8)),
			5948 => std_logic_vector(to_unsigned(78, 8)),
			5949 => std_logic_vector(to_unsigned(69, 8)),
			5950 => std_logic_vector(to_unsigned(91, 8)),
			5951 => std_logic_vector(to_unsigned(222, 8)),
			5952 => std_logic_vector(to_unsigned(55, 8)),
			5953 => std_logic_vector(to_unsigned(79, 8)),
			5954 => std_logic_vector(to_unsigned(5, 8)),
			5955 => std_logic_vector(to_unsigned(162, 8)),
			5956 => std_logic_vector(to_unsigned(19, 8)),
			5957 => std_logic_vector(to_unsigned(122, 8)),
			5958 => std_logic_vector(to_unsigned(109, 8)),
			5959 => std_logic_vector(to_unsigned(15, 8)),
			5960 => std_logic_vector(to_unsigned(38, 8)),
			5961 => std_logic_vector(to_unsigned(10, 8)),
			5962 => std_logic_vector(to_unsigned(252, 8)),
			5963 => std_logic_vector(to_unsigned(136, 8)),
			5964 => std_logic_vector(to_unsigned(149, 8)),
			5965 => std_logic_vector(to_unsigned(168, 8)),
			5966 => std_logic_vector(to_unsigned(168, 8)),
			5967 => std_logic_vector(to_unsigned(130, 8)),
			5968 => std_logic_vector(to_unsigned(12, 8)),
			5969 => std_logic_vector(to_unsigned(27, 8)),
			5970 => std_logic_vector(to_unsigned(252, 8)),
			5971 => std_logic_vector(to_unsigned(149, 8)),
			5972 => std_logic_vector(to_unsigned(162, 8)),
			5973 => std_logic_vector(to_unsigned(109, 8)),
			5974 => std_logic_vector(to_unsigned(48, 8)),
			5975 => std_logic_vector(to_unsigned(202, 8)),
			5976 => std_logic_vector(to_unsigned(151, 8)),
			5977 => std_logic_vector(to_unsigned(131, 8)),
			5978 => std_logic_vector(to_unsigned(154, 8)),
			5979 => std_logic_vector(to_unsigned(148, 8)),
			5980 => std_logic_vector(to_unsigned(243, 8)),
			5981 => std_logic_vector(to_unsigned(186, 8)),
			5982 => std_logic_vector(to_unsigned(251, 8)),
			5983 => std_logic_vector(to_unsigned(110, 8)),
			5984 => std_logic_vector(to_unsigned(189, 8)),
			5985 => std_logic_vector(to_unsigned(78, 8)),
			5986 => std_logic_vector(to_unsigned(151, 8)),
			5987 => std_logic_vector(to_unsigned(162, 8)),
			5988 => std_logic_vector(to_unsigned(6, 8)),
			5989 => std_logic_vector(to_unsigned(123, 8)),
			5990 => std_logic_vector(to_unsigned(170, 8)),
			5991 => std_logic_vector(to_unsigned(60, 8)),
			5992 => std_logic_vector(to_unsigned(10, 8)),
			5993 => std_logic_vector(to_unsigned(5, 8)),
			5994 => std_logic_vector(to_unsigned(215, 8)),
			5995 => std_logic_vector(to_unsigned(187, 8)),
			5996 => std_logic_vector(to_unsigned(158, 8)),
			5997 => std_logic_vector(to_unsigned(150, 8)),
			5998 => std_logic_vector(to_unsigned(2, 8)),
			5999 => std_logic_vector(to_unsigned(88, 8)),
			6000 => std_logic_vector(to_unsigned(153, 8)),
			6001 => std_logic_vector(to_unsigned(28, 8)),
			6002 => std_logic_vector(to_unsigned(45, 8)),
			6003 => std_logic_vector(to_unsigned(196, 8)),
			6004 => std_logic_vector(to_unsigned(197, 8)),
			6005 => std_logic_vector(to_unsigned(114, 8)),
			6006 => std_logic_vector(to_unsigned(92, 8)),
			6007 => std_logic_vector(to_unsigned(246, 8)),
			6008 => std_logic_vector(to_unsigned(177, 8)),
			6009 => std_logic_vector(to_unsigned(235, 8)),
			6010 => std_logic_vector(to_unsigned(251, 8)),
			6011 => std_logic_vector(to_unsigned(28, 8)),
			6012 => std_logic_vector(to_unsigned(111, 8)),
			6013 => std_logic_vector(to_unsigned(88, 8)),
			6014 => std_logic_vector(to_unsigned(126, 8)),
			6015 => std_logic_vector(to_unsigned(116, 8)),
			6016 => std_logic_vector(to_unsigned(197, 8)),
			6017 => std_logic_vector(to_unsigned(121, 8)),
			6018 => std_logic_vector(to_unsigned(145, 8)),
			6019 => std_logic_vector(to_unsigned(84, 8)),
			6020 => std_logic_vector(to_unsigned(111, 8)),
			6021 => std_logic_vector(to_unsigned(100, 8)),
			6022 => std_logic_vector(to_unsigned(155, 8)),
			6023 => std_logic_vector(to_unsigned(183, 8)),
			6024 => std_logic_vector(to_unsigned(226, 8)),
			6025 => std_logic_vector(to_unsigned(131, 8)),
			6026 => std_logic_vector(to_unsigned(42, 8)),
			6027 => std_logic_vector(to_unsigned(84, 8)),
			6028 => std_logic_vector(to_unsigned(146, 8)),
			6029 => std_logic_vector(to_unsigned(184, 8)),
			6030 => std_logic_vector(to_unsigned(211, 8)),
			6031 => std_logic_vector(to_unsigned(251, 8)),
			6032 => std_logic_vector(to_unsigned(121, 8)),
			6033 => std_logic_vector(to_unsigned(145, 8)),
			6034 => std_logic_vector(to_unsigned(79, 8)),
			6035 => std_logic_vector(to_unsigned(113, 8)),
			6036 => std_logic_vector(to_unsigned(139, 8)),
			6037 => std_logic_vector(to_unsigned(15, 8)),
			6038 => std_logic_vector(to_unsigned(135, 8)),
			6039 => std_logic_vector(to_unsigned(135, 8)),
			6040 => std_logic_vector(to_unsigned(232, 8)),
			6041 => std_logic_vector(to_unsigned(165, 8)),
			6042 => std_logic_vector(to_unsigned(45, 8)),
			6043 => std_logic_vector(to_unsigned(87, 8)),
			6044 => std_logic_vector(to_unsigned(32, 8)),
			6045 => std_logic_vector(to_unsigned(51, 8)),
			6046 => std_logic_vector(to_unsigned(26, 8)),
			6047 => std_logic_vector(to_unsigned(197, 8)),
			6048 => std_logic_vector(to_unsigned(13, 8)),
			6049 => std_logic_vector(to_unsigned(148, 8)),
			6050 => std_logic_vector(to_unsigned(252, 8)),
			6051 => std_logic_vector(to_unsigned(142, 8)),
			6052 => std_logic_vector(to_unsigned(210, 8)),
			6053 => std_logic_vector(to_unsigned(89, 8)),
			6054 => std_logic_vector(to_unsigned(27, 8)),
			6055 => std_logic_vector(to_unsigned(186, 8)),
			6056 => std_logic_vector(to_unsigned(169, 8)),
			6057 => std_logic_vector(to_unsigned(148, 8)),
			6058 => std_logic_vector(to_unsigned(9, 8)),
			6059 => std_logic_vector(to_unsigned(222, 8)),
			6060 => std_logic_vector(to_unsigned(192, 8)),
			6061 => std_logic_vector(to_unsigned(12, 8)),
			6062 => std_logic_vector(to_unsigned(4, 8)),
			6063 => std_logic_vector(to_unsigned(224, 8)),
			6064 => std_logic_vector(to_unsigned(91, 8)),
			6065 => std_logic_vector(to_unsigned(67, 8)),
			6066 => std_logic_vector(to_unsigned(50, 8)),
			6067 => std_logic_vector(to_unsigned(236, 8)),
			6068 => std_logic_vector(to_unsigned(201, 8)),
			6069 => std_logic_vector(to_unsigned(160, 8)),
			6070 => std_logic_vector(to_unsigned(115, 8)),
			6071 => std_logic_vector(to_unsigned(101, 8)),
			6072 => std_logic_vector(to_unsigned(166, 8)),
			6073 => std_logic_vector(to_unsigned(115, 8)),
			6074 => std_logic_vector(to_unsigned(237, 8)),
			6075 => std_logic_vector(to_unsigned(82, 8)),
			6076 => std_logic_vector(to_unsigned(126, 8)),
			6077 => std_logic_vector(to_unsigned(161, 8)),
			6078 => std_logic_vector(to_unsigned(80, 8)),
			6079 => std_logic_vector(to_unsigned(84, 8)),
			6080 => std_logic_vector(to_unsigned(50, 8)),
			6081 => std_logic_vector(to_unsigned(87, 8)),
			6082 => std_logic_vector(to_unsigned(131, 8)),
			6083 => std_logic_vector(to_unsigned(65, 8)),
			6084 => std_logic_vector(to_unsigned(233, 8)),
			6085 => std_logic_vector(to_unsigned(158, 8)),
			6086 => std_logic_vector(to_unsigned(73, 8)),
			6087 => std_logic_vector(to_unsigned(21, 8)),
			6088 => std_logic_vector(to_unsigned(218, 8)),
			6089 => std_logic_vector(to_unsigned(85, 8)),
			6090 => std_logic_vector(to_unsigned(35, 8)),
			6091 => std_logic_vector(to_unsigned(73, 8)),
			6092 => std_logic_vector(to_unsigned(85, 8)),
			6093 => std_logic_vector(to_unsigned(156, 8)),
			6094 => std_logic_vector(to_unsigned(140, 8)),
			6095 => std_logic_vector(to_unsigned(210, 8)),
			6096 => std_logic_vector(to_unsigned(193, 8)),
			6097 => std_logic_vector(to_unsigned(219, 8)),
			6098 => std_logic_vector(to_unsigned(155, 8)),
			6099 => std_logic_vector(to_unsigned(245, 8)),
			6100 => std_logic_vector(to_unsigned(46, 8)),
			6101 => std_logic_vector(to_unsigned(90, 8)),
			6102 => std_logic_vector(to_unsigned(144, 8)),
			6103 => std_logic_vector(to_unsigned(112, 8)),
			6104 => std_logic_vector(to_unsigned(51, 8)),
			6105 => std_logic_vector(to_unsigned(34, 8)),
			6106 => std_logic_vector(to_unsigned(87, 8)),
			6107 => std_logic_vector(to_unsigned(183, 8)),
			6108 => std_logic_vector(to_unsigned(81, 8)),
			6109 => std_logic_vector(to_unsigned(56, 8)),
			6110 => std_logic_vector(to_unsigned(160, 8)),
			6111 => std_logic_vector(to_unsigned(26, 8)),
			6112 => std_logic_vector(to_unsigned(213, 8)),
			6113 => std_logic_vector(to_unsigned(158, 8)),
			6114 => std_logic_vector(to_unsigned(92, 8)),
			6115 => std_logic_vector(to_unsigned(224, 8)),
			6116 => std_logic_vector(to_unsigned(104, 8)),
			6117 => std_logic_vector(to_unsigned(6, 8)),
			6118 => std_logic_vector(to_unsigned(79, 8)),
			6119 => std_logic_vector(to_unsigned(115, 8)),
			6120 => std_logic_vector(to_unsigned(240, 8)),
			6121 => std_logic_vector(to_unsigned(120, 8)),
			6122 => std_logic_vector(to_unsigned(50, 8)),
			6123 => std_logic_vector(to_unsigned(58, 8)),
			6124 => std_logic_vector(to_unsigned(16, 8)),
			6125 => std_logic_vector(to_unsigned(124, 8)),
			6126 => std_logic_vector(to_unsigned(255, 8)),
			6127 => std_logic_vector(to_unsigned(120, 8)),
			6128 => std_logic_vector(to_unsigned(182, 8)),
			6129 => std_logic_vector(to_unsigned(118, 8)),
			6130 => std_logic_vector(to_unsigned(187, 8)),
			6131 => std_logic_vector(to_unsigned(77, 8)),
			6132 => std_logic_vector(to_unsigned(187, 8)),
			6133 => std_logic_vector(to_unsigned(18, 8)),
			6134 => std_logic_vector(to_unsigned(255, 8)),
			6135 => std_logic_vector(to_unsigned(118, 8)),
			6136 => std_logic_vector(to_unsigned(58, 8)),
			6137 => std_logic_vector(to_unsigned(196, 8)),
			6138 => std_logic_vector(to_unsigned(136, 8)),
			6139 => std_logic_vector(to_unsigned(47, 8)),
			6140 => std_logic_vector(to_unsigned(218, 8)),
			6141 => std_logic_vector(to_unsigned(234, 8)),
			6142 => std_logic_vector(to_unsigned(171, 8)),
			6143 => std_logic_vector(to_unsigned(171, 8)),
			6144 => std_logic_vector(to_unsigned(217, 8)),
			6145 => std_logic_vector(to_unsigned(91, 8)),
			6146 => std_logic_vector(to_unsigned(223, 8)),
			6147 => std_logic_vector(to_unsigned(76, 8)),
			6148 => std_logic_vector(to_unsigned(155, 8)),
			6149 => std_logic_vector(to_unsigned(18, 8)),
			6150 => std_logic_vector(to_unsigned(234, 8)),
			6151 => std_logic_vector(to_unsigned(118, 8)),
			6152 => std_logic_vector(to_unsigned(147, 8)),
			6153 => std_logic_vector(to_unsigned(114, 8)),
			6154 => std_logic_vector(to_unsigned(32, 8)),
			6155 => std_logic_vector(to_unsigned(30, 8)),
			6156 => std_logic_vector(to_unsigned(168, 8)),
			6157 => std_logic_vector(to_unsigned(59, 8)),
			6158 => std_logic_vector(to_unsigned(70, 8)),
			6159 => std_logic_vector(to_unsigned(107, 8)),
			6160 => std_logic_vector(to_unsigned(220, 8)),
			6161 => std_logic_vector(to_unsigned(186, 8)),
			6162 => std_logic_vector(to_unsigned(137, 8)),
			6163 => std_logic_vector(to_unsigned(139, 8)),
			6164 => std_logic_vector(to_unsigned(192, 8)),
			6165 => std_logic_vector(to_unsigned(26, 8)),
			6166 => std_logic_vector(to_unsigned(90, 8)),
			6167 => std_logic_vector(to_unsigned(213, 8)),
			6168 => std_logic_vector(to_unsigned(127, 8)),
			6169 => std_logic_vector(to_unsigned(235, 8)),
			6170 => std_logic_vector(to_unsigned(3, 8)),
			6171 => std_logic_vector(to_unsigned(93, 8)),
			6172 => std_logic_vector(to_unsigned(45, 8)),
			6173 => std_logic_vector(to_unsigned(187, 8)),
			6174 => std_logic_vector(to_unsigned(111, 8)),
			6175 => std_logic_vector(to_unsigned(216, 8)),
			6176 => std_logic_vector(to_unsigned(82, 8)),
			6177 => std_logic_vector(to_unsigned(9, 8)),
			6178 => std_logic_vector(to_unsigned(212, 8)),
			6179 => std_logic_vector(to_unsigned(111, 8)),
			6180 => std_logic_vector(to_unsigned(248, 8)),
			6181 => std_logic_vector(to_unsigned(237, 8)),
			6182 => std_logic_vector(to_unsigned(7, 8)),
			6183 => std_logic_vector(to_unsigned(156, 8)),
			6184 => std_logic_vector(to_unsigned(84, 8)),
			6185 => std_logic_vector(to_unsigned(249, 8)),
			6186 => std_logic_vector(to_unsigned(203, 8)),
			6187 => std_logic_vector(to_unsigned(0, 8)),
			6188 => std_logic_vector(to_unsigned(223, 8)),
			6189 => std_logic_vector(to_unsigned(2, 8)),
			6190 => std_logic_vector(to_unsigned(240, 8)),
			6191 => std_logic_vector(to_unsigned(185, 8)),
			6192 => std_logic_vector(to_unsigned(112, 8)),
			6193 => std_logic_vector(to_unsigned(122, 8)),
			6194 => std_logic_vector(to_unsigned(88, 8)),
			6195 => std_logic_vector(to_unsigned(95, 8)),
			6196 => std_logic_vector(to_unsigned(214, 8)),
			6197 => std_logic_vector(to_unsigned(219, 8)),
			6198 => std_logic_vector(to_unsigned(75, 8)),
			6199 => std_logic_vector(to_unsigned(211, 8)),
			6200 => std_logic_vector(to_unsigned(125, 8)),
			6201 => std_logic_vector(to_unsigned(59, 8)),
			6202 => std_logic_vector(to_unsigned(172, 8)),
			6203 => std_logic_vector(to_unsigned(68, 8)),
			6204 => std_logic_vector(to_unsigned(36, 8)),
			6205 => std_logic_vector(to_unsigned(65, 8)),
			6206 => std_logic_vector(to_unsigned(199, 8)),
			6207 => std_logic_vector(to_unsigned(111, 8)),
			6208 => std_logic_vector(to_unsigned(205, 8)),
			6209 => std_logic_vector(to_unsigned(115, 8)),
			6210 => std_logic_vector(to_unsigned(103, 8)),
			6211 => std_logic_vector(to_unsigned(121, 8)),
			6212 => std_logic_vector(to_unsigned(151, 8)),
			6213 => std_logic_vector(to_unsigned(246, 8)),
			6214 => std_logic_vector(to_unsigned(47, 8)),
			6215 => std_logic_vector(to_unsigned(96, 8)),
			6216 => std_logic_vector(to_unsigned(104, 8)),
			6217 => std_logic_vector(to_unsigned(164, 8)),
			6218 => std_logic_vector(to_unsigned(73, 8)),
			6219 => std_logic_vector(to_unsigned(122, 8)),
			6220 => std_logic_vector(to_unsigned(57, 8)),
			6221 => std_logic_vector(to_unsigned(48, 8)),
			6222 => std_logic_vector(to_unsigned(12, 8)),
			6223 => std_logic_vector(to_unsigned(246, 8)),
			6224 => std_logic_vector(to_unsigned(88, 8)),
			6225 => std_logic_vector(to_unsigned(15, 8)),
			6226 => std_logic_vector(to_unsigned(38, 8)),
			6227 => std_logic_vector(to_unsigned(34, 8)),
			6228 => std_logic_vector(to_unsigned(52, 8)),
			6229 => std_logic_vector(to_unsigned(106, 8)),
			6230 => std_logic_vector(to_unsigned(199, 8)),
			6231 => std_logic_vector(to_unsigned(2, 8)),
			6232 => std_logic_vector(to_unsigned(145, 8)),
			6233 => std_logic_vector(to_unsigned(41, 8)),
			6234 => std_logic_vector(to_unsigned(72, 8)),
			6235 => std_logic_vector(to_unsigned(64, 8)),
			6236 => std_logic_vector(to_unsigned(40, 8)),
			6237 => std_logic_vector(to_unsigned(14, 8)),
			6238 => std_logic_vector(to_unsigned(249, 8)),
			6239 => std_logic_vector(to_unsigned(45, 8)),
			6240 => std_logic_vector(to_unsigned(212, 8)),
			6241 => std_logic_vector(to_unsigned(49, 8)),
			6242 => std_logic_vector(to_unsigned(81, 8)),
			6243 => std_logic_vector(to_unsigned(0, 8)),
			6244 => std_logic_vector(to_unsigned(161, 8)),
			6245 => std_logic_vector(to_unsigned(70, 8)),
			6246 => std_logic_vector(to_unsigned(58, 8)),
			6247 => std_logic_vector(to_unsigned(206, 8)),
			6248 => std_logic_vector(to_unsigned(181, 8)),
			6249 => std_logic_vector(to_unsigned(59, 8)),
			6250 => std_logic_vector(to_unsigned(171, 8)),
			6251 => std_logic_vector(to_unsigned(105, 8)),
			6252 => std_logic_vector(to_unsigned(4, 8)),
			6253 => std_logic_vector(to_unsigned(173, 8)),
			6254 => std_logic_vector(to_unsigned(123, 8)),
			6255 => std_logic_vector(to_unsigned(231, 8)),
			6256 => std_logic_vector(to_unsigned(23, 8)),
			6257 => std_logic_vector(to_unsigned(254, 8)),
			6258 => std_logic_vector(to_unsigned(53, 8)),
			6259 => std_logic_vector(to_unsigned(180, 8)),
			6260 => std_logic_vector(to_unsigned(247, 8)),
			6261 => std_logic_vector(to_unsigned(3, 8)),
			6262 => std_logic_vector(to_unsigned(87, 8)),
			6263 => std_logic_vector(to_unsigned(89, 8)),
			6264 => std_logic_vector(to_unsigned(103, 8)),
			6265 => std_logic_vector(to_unsigned(47, 8)),
			6266 => std_logic_vector(to_unsigned(85, 8)),
			6267 => std_logic_vector(to_unsigned(69, 8)),
			6268 => std_logic_vector(to_unsigned(231, 8)),
			6269 => std_logic_vector(to_unsigned(211, 8)),
			6270 => std_logic_vector(to_unsigned(231, 8)),
			6271 => std_logic_vector(to_unsigned(175, 8)),
			6272 => std_logic_vector(to_unsigned(184, 8)),
			6273 => std_logic_vector(to_unsigned(6, 8)),
			6274 => std_logic_vector(to_unsigned(95, 8)),
			6275 => std_logic_vector(to_unsigned(18, 8)),
			6276 => std_logic_vector(to_unsigned(96, 8)),
			6277 => std_logic_vector(to_unsigned(151, 8)),
			6278 => std_logic_vector(to_unsigned(209, 8)),
			6279 => std_logic_vector(to_unsigned(198, 8)),
			6280 => std_logic_vector(to_unsigned(176, 8)),
			6281 => std_logic_vector(to_unsigned(141, 8)),
			6282 => std_logic_vector(to_unsigned(171, 8)),
			6283 => std_logic_vector(to_unsigned(186, 8)),
			6284 => std_logic_vector(to_unsigned(195, 8)),
			6285 => std_logic_vector(to_unsigned(53, 8)),
			6286 => std_logic_vector(to_unsigned(46, 8)),
			6287 => std_logic_vector(to_unsigned(123, 8)),
			6288 => std_logic_vector(to_unsigned(247, 8)),
			6289 => std_logic_vector(to_unsigned(36, 8)),
			6290 => std_logic_vector(to_unsigned(108, 8)),
			6291 => std_logic_vector(to_unsigned(162, 8)),
			6292 => std_logic_vector(to_unsigned(111, 8)),
			6293 => std_logic_vector(to_unsigned(32, 8)),
			6294 => std_logic_vector(to_unsigned(141, 8)),
			6295 => std_logic_vector(to_unsigned(50, 8)),
			6296 => std_logic_vector(to_unsigned(169, 8)),
			6297 => std_logic_vector(to_unsigned(203, 8)),
			6298 => std_logic_vector(to_unsigned(215, 8)),
			6299 => std_logic_vector(to_unsigned(209, 8)),
			6300 => std_logic_vector(to_unsigned(167, 8)),
			6301 => std_logic_vector(to_unsigned(209, 8)),
			6302 => std_logic_vector(to_unsigned(119, 8)),
			6303 => std_logic_vector(to_unsigned(69, 8)),
			6304 => std_logic_vector(to_unsigned(180, 8)),
			6305 => std_logic_vector(to_unsigned(33, 8)),
			6306 => std_logic_vector(to_unsigned(170, 8)),
			6307 => std_logic_vector(to_unsigned(206, 8)),
			6308 => std_logic_vector(to_unsigned(213, 8)),
			6309 => std_logic_vector(to_unsigned(115, 8)),
			6310 => std_logic_vector(to_unsigned(60, 8)),
			6311 => std_logic_vector(to_unsigned(193, 8)),
			6312 => std_logic_vector(to_unsigned(244, 8)),
			6313 => std_logic_vector(to_unsigned(109, 8)),
			6314 => std_logic_vector(to_unsigned(187, 8)),
			6315 => std_logic_vector(to_unsigned(200, 8)),
			6316 => std_logic_vector(to_unsigned(162, 8)),
			6317 => std_logic_vector(to_unsigned(200, 8)),
			6318 => std_logic_vector(to_unsigned(33, 8)),
			6319 => std_logic_vector(to_unsigned(58, 8)),
			6320 => std_logic_vector(to_unsigned(25, 8)),
			6321 => std_logic_vector(to_unsigned(226, 8)),
			6322 => std_logic_vector(to_unsigned(112, 8)),
			6323 => std_logic_vector(to_unsigned(141, 8)),
			6324 => std_logic_vector(to_unsigned(210, 8)),
			6325 => std_logic_vector(to_unsigned(49, 8)),
			6326 => std_logic_vector(to_unsigned(163, 8)),
			6327 => std_logic_vector(to_unsigned(1, 8)),
			6328 => std_logic_vector(to_unsigned(138, 8)),
			6329 => std_logic_vector(to_unsigned(214, 8)),
			6330 => std_logic_vector(to_unsigned(61, 8)),
			6331 => std_logic_vector(to_unsigned(45, 8)),
			6332 => std_logic_vector(to_unsigned(218, 8)),
			6333 => std_logic_vector(to_unsigned(240, 8)),
			6334 => std_logic_vector(to_unsigned(56, 8)),
			6335 => std_logic_vector(to_unsigned(157, 8)),
			6336 => std_logic_vector(to_unsigned(151, 8)),
			6337 => std_logic_vector(to_unsigned(93, 8)),
			6338 => std_logic_vector(to_unsigned(85, 8)),
			6339 => std_logic_vector(to_unsigned(244, 8)),
			6340 => std_logic_vector(to_unsigned(221, 8)),
			6341 => std_logic_vector(to_unsigned(218, 8)),
			6342 => std_logic_vector(to_unsigned(245, 8)),
			6343 => std_logic_vector(to_unsigned(250, 8)),
			6344 => std_logic_vector(to_unsigned(178, 8)),
			6345 => std_logic_vector(to_unsigned(199, 8)),
			6346 => std_logic_vector(to_unsigned(128, 8)),
			6347 => std_logic_vector(to_unsigned(168, 8)),
			6348 => std_logic_vector(to_unsigned(29, 8)),
			6349 => std_logic_vector(to_unsigned(185, 8)),
			6350 => std_logic_vector(to_unsigned(102, 8)),
			6351 => std_logic_vector(to_unsigned(50, 8)),
			6352 => std_logic_vector(to_unsigned(235, 8)),
			6353 => std_logic_vector(to_unsigned(77, 8)),
			6354 => std_logic_vector(to_unsigned(224, 8)),
			6355 => std_logic_vector(to_unsigned(82, 8)),
			6356 => std_logic_vector(to_unsigned(22, 8)),
			6357 => std_logic_vector(to_unsigned(3, 8)),
			6358 => std_logic_vector(to_unsigned(148, 8)),
			6359 => std_logic_vector(to_unsigned(35, 8)),
			6360 => std_logic_vector(to_unsigned(22, 8)),
			6361 => std_logic_vector(to_unsigned(196, 8)),
			6362 => std_logic_vector(to_unsigned(18, 8)),
			6363 => std_logic_vector(to_unsigned(41, 8)),
			6364 => std_logic_vector(to_unsigned(236, 8)),
			6365 => std_logic_vector(to_unsigned(164, 8)),
			6366 => std_logic_vector(to_unsigned(162, 8)),
			6367 => std_logic_vector(to_unsigned(248, 8)),
			6368 => std_logic_vector(to_unsigned(161, 8)),
			6369 => std_logic_vector(to_unsigned(200, 8)),
			6370 => std_logic_vector(to_unsigned(2, 8)),
			6371 => std_logic_vector(to_unsigned(218, 8)),
			6372 => std_logic_vector(to_unsigned(142, 8)),
			6373 => std_logic_vector(to_unsigned(177, 8)),
			6374 => std_logic_vector(to_unsigned(161, 8)),
			6375 => std_logic_vector(to_unsigned(186, 8)),
			6376 => std_logic_vector(to_unsigned(184, 8)),
			6377 => std_logic_vector(to_unsigned(24, 8)),
			6378 => std_logic_vector(to_unsigned(53, 8)),
			6379 => std_logic_vector(to_unsigned(232, 8)),
			6380 => std_logic_vector(to_unsigned(151, 8)),
			6381 => std_logic_vector(to_unsigned(247, 8)),
			6382 => std_logic_vector(to_unsigned(44, 8)),
			6383 => std_logic_vector(to_unsigned(137, 8)),
			6384 => std_logic_vector(to_unsigned(119, 8)),
			6385 => std_logic_vector(to_unsigned(185, 8)),
			6386 => std_logic_vector(to_unsigned(250, 8)),
			6387 => std_logic_vector(to_unsigned(99, 8)),
			6388 => std_logic_vector(to_unsigned(60, 8)),
			6389 => std_logic_vector(to_unsigned(206, 8)),
			6390 => std_logic_vector(to_unsigned(53, 8)),
			6391 => std_logic_vector(to_unsigned(176, 8)),
			6392 => std_logic_vector(to_unsigned(20, 8)),
			6393 => std_logic_vector(to_unsigned(226, 8)),
			6394 => std_logic_vector(to_unsigned(255, 8)),
			6395 => std_logic_vector(to_unsigned(191, 8)),
			6396 => std_logic_vector(to_unsigned(244, 8)),
			6397 => std_logic_vector(to_unsigned(178, 8)),
			6398 => std_logic_vector(to_unsigned(49, 8)),
			6399 => std_logic_vector(to_unsigned(238, 8)),
			6400 => std_logic_vector(to_unsigned(145, 8)),
			6401 => std_logic_vector(to_unsigned(91, 8)),
			6402 => std_logic_vector(to_unsigned(144, 8)),
			6403 => std_logic_vector(to_unsigned(160, 8)),
			6404 => std_logic_vector(to_unsigned(68, 8)),
			6405 => std_logic_vector(to_unsigned(131, 8)),
			6406 => std_logic_vector(to_unsigned(164, 8)),
			6407 => std_logic_vector(to_unsigned(38, 8)),
			6408 => std_logic_vector(to_unsigned(88, 8)),
			6409 => std_logic_vector(to_unsigned(213, 8)),
			6410 => std_logic_vector(to_unsigned(78, 8)),
			6411 => std_logic_vector(to_unsigned(25, 8)),
			6412 => std_logic_vector(to_unsigned(180, 8)),
			6413 => std_logic_vector(to_unsigned(186, 8)),
			6414 => std_logic_vector(to_unsigned(174, 8)),
			6415 => std_logic_vector(to_unsigned(12, 8)),
			6416 => std_logic_vector(to_unsigned(150, 8)),
			6417 => std_logic_vector(to_unsigned(83, 8)),
			6418 => std_logic_vector(to_unsigned(154, 8)),
			6419 => std_logic_vector(to_unsigned(83, 8)),
			6420 => std_logic_vector(to_unsigned(105, 8)),
			6421 => std_logic_vector(to_unsigned(255, 8)),
			6422 => std_logic_vector(to_unsigned(238, 8)),
			6423 => std_logic_vector(to_unsigned(204, 8)),
			6424 => std_logic_vector(to_unsigned(39, 8)),
			6425 => std_logic_vector(to_unsigned(71, 8)),
			6426 => std_logic_vector(to_unsigned(191, 8)),
			6427 => std_logic_vector(to_unsigned(196, 8)),
			6428 => std_logic_vector(to_unsigned(48, 8)),
			6429 => std_logic_vector(to_unsigned(25, 8)),
			6430 => std_logic_vector(to_unsigned(208, 8)),
			6431 => std_logic_vector(to_unsigned(8, 8)),
			6432 => std_logic_vector(to_unsigned(225, 8)),
			6433 => std_logic_vector(to_unsigned(231, 8)),
			6434 => std_logic_vector(to_unsigned(195, 8)),
			6435 => std_logic_vector(to_unsigned(28, 8)),
			6436 => std_logic_vector(to_unsigned(153, 8)),
			6437 => std_logic_vector(to_unsigned(129, 8)),
			6438 => std_logic_vector(to_unsigned(195, 8)),
			6439 => std_logic_vector(to_unsigned(133, 8)),
			6440 => std_logic_vector(to_unsigned(75, 8)),
			6441 => std_logic_vector(to_unsigned(90, 8)),
			6442 => std_logic_vector(to_unsigned(116, 8)),
			6443 => std_logic_vector(to_unsigned(133, 8)),
			6444 => std_logic_vector(to_unsigned(215, 8)),
			6445 => std_logic_vector(to_unsigned(211, 8)),
			6446 => std_logic_vector(to_unsigned(60, 8)),
			6447 => std_logic_vector(to_unsigned(228, 8)),
			6448 => std_logic_vector(to_unsigned(83, 8)),
			6449 => std_logic_vector(to_unsigned(50, 8)),
			6450 => std_logic_vector(to_unsigned(6, 8)),
			6451 => std_logic_vector(to_unsigned(66, 8)),
			6452 => std_logic_vector(to_unsigned(160, 8)),
			6453 => std_logic_vector(to_unsigned(178, 8)),
			6454 => std_logic_vector(to_unsigned(139, 8)),
			6455 => std_logic_vector(to_unsigned(2, 8)),
			6456 => std_logic_vector(to_unsigned(222, 8)),
			6457 => std_logic_vector(to_unsigned(111, 8)),
			6458 => std_logic_vector(to_unsigned(144, 8)),
			6459 => std_logic_vector(to_unsigned(173, 8)),
			6460 => std_logic_vector(to_unsigned(101, 8)),
			6461 => std_logic_vector(to_unsigned(246, 8)),
			6462 => std_logic_vector(to_unsigned(255, 8)),
			6463 => std_logic_vector(to_unsigned(148, 8)),
			6464 => std_logic_vector(to_unsigned(47, 8)),
			6465 => std_logic_vector(to_unsigned(1, 8)),
			6466 => std_logic_vector(to_unsigned(50, 8)),
			6467 => std_logic_vector(to_unsigned(120, 8)),
			6468 => std_logic_vector(to_unsigned(71, 8)),
			6469 => std_logic_vector(to_unsigned(56, 8)),
			6470 => std_logic_vector(to_unsigned(97, 8)),
			6471 => std_logic_vector(to_unsigned(234, 8)),
			6472 => std_logic_vector(to_unsigned(126, 8)),
			6473 => std_logic_vector(to_unsigned(76, 8)),
			6474 => std_logic_vector(to_unsigned(192, 8)),
			6475 => std_logic_vector(to_unsigned(124, 8)),
			6476 => std_logic_vector(to_unsigned(50, 8)),
			6477 => std_logic_vector(to_unsigned(120, 8)),
			6478 => std_logic_vector(to_unsigned(41, 8)),
			6479 => std_logic_vector(to_unsigned(217, 8)),
			6480 => std_logic_vector(to_unsigned(243, 8)),
			6481 => std_logic_vector(to_unsigned(208, 8)),
			6482 => std_logic_vector(to_unsigned(243, 8)),
			6483 => std_logic_vector(to_unsigned(58, 8)),
			6484 => std_logic_vector(to_unsigned(116, 8)),
			6485 => std_logic_vector(to_unsigned(248, 8)),
			6486 => std_logic_vector(to_unsigned(64, 8)),
			6487 => std_logic_vector(to_unsigned(175, 8)),
			6488 => std_logic_vector(to_unsigned(249, 8)),
			6489 => std_logic_vector(to_unsigned(76, 8)),
			6490 => std_logic_vector(to_unsigned(12, 8)),
			6491 => std_logic_vector(to_unsigned(234, 8)),
			6492 => std_logic_vector(to_unsigned(173, 8)),
			6493 => std_logic_vector(to_unsigned(183, 8)),
			6494 => std_logic_vector(to_unsigned(194, 8)),
			6495 => std_logic_vector(to_unsigned(178, 8)),
			6496 => std_logic_vector(to_unsigned(0, 8)),
			6497 => std_logic_vector(to_unsigned(36, 8)),
			6498 => std_logic_vector(to_unsigned(145, 8)),
			6499 => std_logic_vector(to_unsigned(119, 8)),
			6500 => std_logic_vector(to_unsigned(229, 8)),
			6501 => std_logic_vector(to_unsigned(58, 8)),
			6502 => std_logic_vector(to_unsigned(119, 8)),
			6503 => std_logic_vector(to_unsigned(200, 8)),
			6504 => std_logic_vector(to_unsigned(124, 8)),
			6505 => std_logic_vector(to_unsigned(146, 8)),
			6506 => std_logic_vector(to_unsigned(51, 8)),
			6507 => std_logic_vector(to_unsigned(148, 8)),
			6508 => std_logic_vector(to_unsigned(21, 8)),
			6509 => std_logic_vector(to_unsigned(90, 8)),
			6510 => std_logic_vector(to_unsigned(249, 8)),
			6511 => std_logic_vector(to_unsigned(217, 8)),
			6512 => std_logic_vector(to_unsigned(137, 8)),
			6513 => std_logic_vector(to_unsigned(163, 8)),
			6514 => std_logic_vector(to_unsigned(17, 8)),
			6515 => std_logic_vector(to_unsigned(226, 8)),
			6516 => std_logic_vector(to_unsigned(180, 8)),
			6517 => std_logic_vector(to_unsigned(165, 8)),
			6518 => std_logic_vector(to_unsigned(7, 8)),
			6519 => std_logic_vector(to_unsigned(233, 8)),
			6520 => std_logic_vector(to_unsigned(235, 8)),
			6521 => std_logic_vector(to_unsigned(28, 8)),
			6522 => std_logic_vector(to_unsigned(27, 8)),
			6523 => std_logic_vector(to_unsigned(65, 8)),
			6524 => std_logic_vector(to_unsigned(11, 8)),
			6525 => std_logic_vector(to_unsigned(183, 8)),
			6526 => std_logic_vector(to_unsigned(250, 8)),
			6527 => std_logic_vector(to_unsigned(75, 8)),
			6528 => std_logic_vector(to_unsigned(159, 8)),
			6529 => std_logic_vector(to_unsigned(247, 8)),
			6530 => std_logic_vector(to_unsigned(196, 8)),
			6531 => std_logic_vector(to_unsigned(206, 8)),
			6532 => std_logic_vector(to_unsigned(249, 8)),
			6533 => std_logic_vector(to_unsigned(134, 8)),
			6534 => std_logic_vector(to_unsigned(153, 8)),
			6535 => std_logic_vector(to_unsigned(75, 8)),
			6536 => std_logic_vector(to_unsigned(130, 8)),
			6537 => std_logic_vector(to_unsigned(8, 8)),
			6538 => std_logic_vector(to_unsigned(119, 8)),
			6539 => std_logic_vector(to_unsigned(48, 8)),
			6540 => std_logic_vector(to_unsigned(73, 8)),
			6541 => std_logic_vector(to_unsigned(149, 8)),
			6542 => std_logic_vector(to_unsigned(196, 8)),
			6543 => std_logic_vector(to_unsigned(148, 8)),
			6544 => std_logic_vector(to_unsigned(245, 8)),
			6545 => std_logic_vector(to_unsigned(96, 8)),
			6546 => std_logic_vector(to_unsigned(133, 8)),
			6547 => std_logic_vector(to_unsigned(207, 8)),
			6548 => std_logic_vector(to_unsigned(180, 8)),
			6549 => std_logic_vector(to_unsigned(85, 8)),
			6550 => std_logic_vector(to_unsigned(136, 8)),
			6551 => std_logic_vector(to_unsigned(164, 8)),
			6552 => std_logic_vector(to_unsigned(229, 8)),
			6553 => std_logic_vector(to_unsigned(139, 8)),
			6554 => std_logic_vector(to_unsigned(29, 8)),
			6555 => std_logic_vector(to_unsigned(30, 8)),
			6556 => std_logic_vector(to_unsigned(40, 8)),
			6557 => std_logic_vector(to_unsigned(174, 8)),
			6558 => std_logic_vector(to_unsigned(152, 8)),
			6559 => std_logic_vector(to_unsigned(77, 8)),
			6560 => std_logic_vector(to_unsigned(153, 8)),
			6561 => std_logic_vector(to_unsigned(44, 8)),
			6562 => std_logic_vector(to_unsigned(178, 8)),
			6563 => std_logic_vector(to_unsigned(155, 8)),
			6564 => std_logic_vector(to_unsigned(29, 8)),
			6565 => std_logic_vector(to_unsigned(116, 8)),
			6566 => std_logic_vector(to_unsigned(212, 8)),
			6567 => std_logic_vector(to_unsigned(75, 8)),
			6568 => std_logic_vector(to_unsigned(34, 8)),
			6569 => std_logic_vector(to_unsigned(217, 8)),
			6570 => std_logic_vector(to_unsigned(241, 8)),
			6571 => std_logic_vector(to_unsigned(105, 8)),
			6572 => std_logic_vector(to_unsigned(181, 8)),
			6573 => std_logic_vector(to_unsigned(66, 8)),
			6574 => std_logic_vector(to_unsigned(56, 8)),
			6575 => std_logic_vector(to_unsigned(160, 8)),
			6576 => std_logic_vector(to_unsigned(158, 8)),
			6577 => std_logic_vector(to_unsigned(217, 8)),
			6578 => std_logic_vector(to_unsigned(255, 8)),
			6579 => std_logic_vector(to_unsigned(252, 8)),
			6580 => std_logic_vector(to_unsigned(111, 8)),
			6581 => std_logic_vector(to_unsigned(43, 8)),
			6582 => std_logic_vector(to_unsigned(127, 8)),
			6583 => std_logic_vector(to_unsigned(223, 8)),
			6584 => std_logic_vector(to_unsigned(17, 8)),
			6585 => std_logic_vector(to_unsigned(145, 8)),
			6586 => std_logic_vector(to_unsigned(178, 8)),
			6587 => std_logic_vector(to_unsigned(18, 8)),
			6588 => std_logic_vector(to_unsigned(244, 8)),
			6589 => std_logic_vector(to_unsigned(177, 8)),
			6590 => std_logic_vector(to_unsigned(77, 8)),
			6591 => std_logic_vector(to_unsigned(76, 8)),
			6592 => std_logic_vector(to_unsigned(227, 8)),
			6593 => std_logic_vector(to_unsigned(2, 8)),
			6594 => std_logic_vector(to_unsigned(10, 8)),
			6595 => std_logic_vector(to_unsigned(209, 8)),
			6596 => std_logic_vector(to_unsigned(209, 8)),
			6597 => std_logic_vector(to_unsigned(206, 8)),
			6598 => std_logic_vector(to_unsigned(89, 8)),
			6599 => std_logic_vector(to_unsigned(60, 8)),
			6600 => std_logic_vector(to_unsigned(61, 8)),
			6601 => std_logic_vector(to_unsigned(111, 8)),
			6602 => std_logic_vector(to_unsigned(184, 8)),
			6603 => std_logic_vector(to_unsigned(212, 8)),
			6604 => std_logic_vector(to_unsigned(13, 8)),
			6605 => std_logic_vector(to_unsigned(231, 8)),
			6606 => std_logic_vector(to_unsigned(66, 8)),
			6607 => std_logic_vector(to_unsigned(228, 8)),
			6608 => std_logic_vector(to_unsigned(196, 8)),
			6609 => std_logic_vector(to_unsigned(33, 8)),
			6610 => std_logic_vector(to_unsigned(208, 8)),
			6611 => std_logic_vector(to_unsigned(146, 8)),
			6612 => std_logic_vector(to_unsigned(52, 8)),
			6613 => std_logic_vector(to_unsigned(208, 8)),
			6614 => std_logic_vector(to_unsigned(169, 8)),
			6615 => std_logic_vector(to_unsigned(93, 8)),
			6616 => std_logic_vector(to_unsigned(233, 8)),
			6617 => std_logic_vector(to_unsigned(248, 8)),
			6618 => std_logic_vector(to_unsigned(34, 8)),
			6619 => std_logic_vector(to_unsigned(144, 8)),
			6620 => std_logic_vector(to_unsigned(246, 8)),
			6621 => std_logic_vector(to_unsigned(150, 8)),
			6622 => std_logic_vector(to_unsigned(111, 8)),
			6623 => std_logic_vector(to_unsigned(233, 8)),
			6624 => std_logic_vector(to_unsigned(121, 8)),
			6625 => std_logic_vector(to_unsigned(40, 8)),
			6626 => std_logic_vector(to_unsigned(251, 8)),
			6627 => std_logic_vector(to_unsigned(22, 8)),
			6628 => std_logic_vector(to_unsigned(4, 8)),
			6629 => std_logic_vector(to_unsigned(65, 8)),
			6630 => std_logic_vector(to_unsigned(104, 8)),
			6631 => std_logic_vector(to_unsigned(61, 8)),
			6632 => std_logic_vector(to_unsigned(101, 8)),
			6633 => std_logic_vector(to_unsigned(166, 8)),
			6634 => std_logic_vector(to_unsigned(43, 8)),
			6635 => std_logic_vector(to_unsigned(117, 8)),
			6636 => std_logic_vector(to_unsigned(218, 8)),
			6637 => std_logic_vector(to_unsigned(215, 8)),
			6638 => std_logic_vector(to_unsigned(82, 8)),
			6639 => std_logic_vector(to_unsigned(81, 8)),
			6640 => std_logic_vector(to_unsigned(6, 8)),
			6641 => std_logic_vector(to_unsigned(30, 8)),
			6642 => std_logic_vector(to_unsigned(245, 8)),
			6643 => std_logic_vector(to_unsigned(154, 8)),
			6644 => std_logic_vector(to_unsigned(31, 8)),
			6645 => std_logic_vector(to_unsigned(75, 8)),
			6646 => std_logic_vector(to_unsigned(184, 8)),
			6647 => std_logic_vector(to_unsigned(94, 8)),
			6648 => std_logic_vector(to_unsigned(216, 8)),
			6649 => std_logic_vector(to_unsigned(28, 8)),
			6650 => std_logic_vector(to_unsigned(218, 8)),
			6651 => std_logic_vector(to_unsigned(145, 8)),
			6652 => std_logic_vector(to_unsigned(179, 8)),
			6653 => std_logic_vector(to_unsigned(199, 8)),
			6654 => std_logic_vector(to_unsigned(247, 8)),
			6655 => std_logic_vector(to_unsigned(205, 8)),
			6656 => std_logic_vector(to_unsigned(56, 8)),
			6657 => std_logic_vector(to_unsigned(214, 8)),
			6658 => std_logic_vector(to_unsigned(21, 8)),
			6659 => std_logic_vector(to_unsigned(45, 8)),
			6660 => std_logic_vector(to_unsigned(183, 8)),
			6661 => std_logic_vector(to_unsigned(99, 8)),
			6662 => std_logic_vector(to_unsigned(214, 8)),
			6663 => std_logic_vector(to_unsigned(139, 8)),
			6664 => std_logic_vector(to_unsigned(99, 8)),
			6665 => std_logic_vector(to_unsigned(200, 8)),
			6666 => std_logic_vector(to_unsigned(197, 8)),
			6667 => std_logic_vector(to_unsigned(76, 8)),
			6668 => std_logic_vector(to_unsigned(188, 8)),
			6669 => std_logic_vector(to_unsigned(56, 8)),
			6670 => std_logic_vector(to_unsigned(164, 8)),
			6671 => std_logic_vector(to_unsigned(243, 8)),
			6672 => std_logic_vector(to_unsigned(174, 8)),
			6673 => std_logic_vector(to_unsigned(10, 8)),
			6674 => std_logic_vector(to_unsigned(17, 8)),
			6675 => std_logic_vector(to_unsigned(227, 8)),
			6676 => std_logic_vector(to_unsigned(79, 8)),
			6677 => std_logic_vector(to_unsigned(205, 8)),
			6678 => std_logic_vector(to_unsigned(140, 8)),
			6679 => std_logic_vector(to_unsigned(73, 8)),
			6680 => std_logic_vector(to_unsigned(118, 8)),
			6681 => std_logic_vector(to_unsigned(169, 8)),
			6682 => std_logic_vector(to_unsigned(137, 8)),
			6683 => std_logic_vector(to_unsigned(166, 8)),
			6684 => std_logic_vector(to_unsigned(84, 8)),
			6685 => std_logic_vector(to_unsigned(107, 8)),
			6686 => std_logic_vector(to_unsigned(108, 8)),
			6687 => std_logic_vector(to_unsigned(222, 8)),
			6688 => std_logic_vector(to_unsigned(254, 8)),
			6689 => std_logic_vector(to_unsigned(85, 8)),
			6690 => std_logic_vector(to_unsigned(158, 8)),
			6691 => std_logic_vector(to_unsigned(228, 8)),
			6692 => std_logic_vector(to_unsigned(65, 8)),
			6693 => std_logic_vector(to_unsigned(248, 8)),
			6694 => std_logic_vector(to_unsigned(217, 8)),
			6695 => std_logic_vector(to_unsigned(66, 8)),
			6696 => std_logic_vector(to_unsigned(92, 8)),
			6697 => std_logic_vector(to_unsigned(210, 8)),
			6698 => std_logic_vector(to_unsigned(43, 8)),
			6699 => std_logic_vector(to_unsigned(187, 8)),
			6700 => std_logic_vector(to_unsigned(108, 8)),
			6701 => std_logic_vector(to_unsigned(81, 8)),
			6702 => std_logic_vector(to_unsigned(249, 8)),
			6703 => std_logic_vector(to_unsigned(96, 8)),
			6704 => std_logic_vector(to_unsigned(60, 8)),
			6705 => std_logic_vector(to_unsigned(228, 8)),
			6706 => std_logic_vector(to_unsigned(216, 8)),
			6707 => std_logic_vector(to_unsigned(190, 8)),
			6708 => std_logic_vector(to_unsigned(154, 8)),
			6709 => std_logic_vector(to_unsigned(14, 8)),
			6710 => std_logic_vector(to_unsigned(30, 8)),
			6711 => std_logic_vector(to_unsigned(157, 8)),
			6712 => std_logic_vector(to_unsigned(199, 8)),
			6713 => std_logic_vector(to_unsigned(254, 8)),
			6714 => std_logic_vector(to_unsigned(151, 8)),
			6715 => std_logic_vector(to_unsigned(49, 8)),
			6716 => std_logic_vector(to_unsigned(243, 8)),
			6717 => std_logic_vector(to_unsigned(39, 8)),
			6718 => std_logic_vector(to_unsigned(221, 8)),
			6719 => std_logic_vector(to_unsigned(254, 8)),
			6720 => std_logic_vector(to_unsigned(254, 8)),
			6721 => std_logic_vector(to_unsigned(174, 8)),
			6722 => std_logic_vector(to_unsigned(190, 8)),
			6723 => std_logic_vector(to_unsigned(66, 8)),
			6724 => std_logic_vector(to_unsigned(157, 8)),
			6725 => std_logic_vector(to_unsigned(78, 8)),
			6726 => std_logic_vector(to_unsigned(151, 8)),
			6727 => std_logic_vector(to_unsigned(240, 8)),
			6728 => std_logic_vector(to_unsigned(174, 8)),
			6729 => std_logic_vector(to_unsigned(16, 8)),
			6730 => std_logic_vector(to_unsigned(192, 8)),
			6731 => std_logic_vector(to_unsigned(173, 8)),
			6732 => std_logic_vector(to_unsigned(35, 8)),
			6733 => std_logic_vector(to_unsigned(35, 8)),
			6734 => std_logic_vector(to_unsigned(78, 8)),
			6735 => std_logic_vector(to_unsigned(164, 8)),
			6736 => std_logic_vector(to_unsigned(199, 8)),
			6737 => std_logic_vector(to_unsigned(238, 8)),
			6738 => std_logic_vector(to_unsigned(59, 8)),
			6739 => std_logic_vector(to_unsigned(46, 8)),
			6740 => std_logic_vector(to_unsigned(124, 8)),
			6741 => std_logic_vector(to_unsigned(169, 8)),
			6742 => std_logic_vector(to_unsigned(254, 8)),
			6743 => std_logic_vector(to_unsigned(233, 8)),
			6744 => std_logic_vector(to_unsigned(47, 8)),
			6745 => std_logic_vector(to_unsigned(112, 8)),
			6746 => std_logic_vector(to_unsigned(37, 8)),
			6747 => std_logic_vector(to_unsigned(152, 8)),
			6748 => std_logic_vector(to_unsigned(84, 8)),
			6749 => std_logic_vector(to_unsigned(53, 8)),
			6750 => std_logic_vector(to_unsigned(118, 8)),
			6751 => std_logic_vector(to_unsigned(202, 8)),
			6752 => std_logic_vector(to_unsigned(96, 8)),
			6753 => std_logic_vector(to_unsigned(72, 8)),
			6754 => std_logic_vector(to_unsigned(159, 8)),
			6755 => std_logic_vector(to_unsigned(134, 8)),
			6756 => std_logic_vector(to_unsigned(202, 8)),
			6757 => std_logic_vector(to_unsigned(102, 8)),
			6758 => std_logic_vector(to_unsigned(35, 8)),
			6759 => std_logic_vector(to_unsigned(124, 8)),
			6760 => std_logic_vector(to_unsigned(82, 8)),
			6761 => std_logic_vector(to_unsigned(60, 8)),
			6762 => std_logic_vector(to_unsigned(193, 8)),
			6763 => std_logic_vector(to_unsigned(53, 8)),
			6764 => std_logic_vector(to_unsigned(172, 8)),
			6765 => std_logic_vector(to_unsigned(124, 8)),
			6766 => std_logic_vector(to_unsigned(176, 8)),
			6767 => std_logic_vector(to_unsigned(33, 8)),
			6768 => std_logic_vector(to_unsigned(140, 8)),
			6769 => std_logic_vector(to_unsigned(191, 8)),
			6770 => std_logic_vector(to_unsigned(22, 8)),
			6771 => std_logic_vector(to_unsigned(134, 8)),
			6772 => std_logic_vector(to_unsigned(111, 8)),
			6773 => std_logic_vector(to_unsigned(122, 8)),
			6774 => std_logic_vector(to_unsigned(101, 8)),
			6775 => std_logic_vector(to_unsigned(126, 8)),
			6776 => std_logic_vector(to_unsigned(112, 8)),
			6777 => std_logic_vector(to_unsigned(99, 8)),
			6778 => std_logic_vector(to_unsigned(226, 8)),
			6779 => std_logic_vector(to_unsigned(210, 8)),
			6780 => std_logic_vector(to_unsigned(175, 8)),
			6781 => std_logic_vector(to_unsigned(133, 8)),
			6782 => std_logic_vector(to_unsigned(71, 8)),
			6783 => std_logic_vector(to_unsigned(40, 8)),
			6784 => std_logic_vector(to_unsigned(93, 8)),
			6785 => std_logic_vector(to_unsigned(161, 8)),
			6786 => std_logic_vector(to_unsigned(84, 8)),
			6787 => std_logic_vector(to_unsigned(11, 8)),
			6788 => std_logic_vector(to_unsigned(248, 8)),
			6789 => std_logic_vector(to_unsigned(139, 8)),
			6790 => std_logic_vector(to_unsigned(250, 8)),
			6791 => std_logic_vector(to_unsigned(5, 8)),
			6792 => std_logic_vector(to_unsigned(30, 8)),
			6793 => std_logic_vector(to_unsigned(83, 8)),
			6794 => std_logic_vector(to_unsigned(3, 8)),
			6795 => std_logic_vector(to_unsigned(50, 8)),
			6796 => std_logic_vector(to_unsigned(247, 8)),
			6797 => std_logic_vector(to_unsigned(51, 8)),
			6798 => std_logic_vector(to_unsigned(154, 8)),
			6799 => std_logic_vector(to_unsigned(173, 8)),
			6800 => std_logic_vector(to_unsigned(219, 8)),
			6801 => std_logic_vector(to_unsigned(136, 8)),
			6802 => std_logic_vector(to_unsigned(69, 8)),
			6803 => std_logic_vector(to_unsigned(71, 8)),
			6804 => std_logic_vector(to_unsigned(94, 8)),
			6805 => std_logic_vector(to_unsigned(105, 8)),
			6806 => std_logic_vector(to_unsigned(182, 8)),
			6807 => std_logic_vector(to_unsigned(51, 8)),
			6808 => std_logic_vector(to_unsigned(145, 8)),
			6809 => std_logic_vector(to_unsigned(20, 8)),
			6810 => std_logic_vector(to_unsigned(89, 8)),
			6811 => std_logic_vector(to_unsigned(15, 8)),
			6812 => std_logic_vector(to_unsigned(149, 8)),
			6813 => std_logic_vector(to_unsigned(110, 8)),
			6814 => std_logic_vector(to_unsigned(196, 8)),
			6815 => std_logic_vector(to_unsigned(65, 8)),
			6816 => std_logic_vector(to_unsigned(47, 8)),
			6817 => std_logic_vector(to_unsigned(48, 8)),
			6818 => std_logic_vector(to_unsigned(77, 8)),
			6819 => std_logic_vector(to_unsigned(153, 8)),
			6820 => std_logic_vector(to_unsigned(190, 8)),
			6821 => std_logic_vector(to_unsigned(243, 8)),
			6822 => std_logic_vector(to_unsigned(177, 8)),
			6823 => std_logic_vector(to_unsigned(240, 8)),
			6824 => std_logic_vector(to_unsigned(120, 8)),
			6825 => std_logic_vector(to_unsigned(66, 8)),
			6826 => std_logic_vector(to_unsigned(249, 8)),
			6827 => std_logic_vector(to_unsigned(169, 8)),
			6828 => std_logic_vector(to_unsigned(193, 8)),
			6829 => std_logic_vector(to_unsigned(37, 8)),
			6830 => std_logic_vector(to_unsigned(228, 8)),
			6831 => std_logic_vector(to_unsigned(121, 8)),
			6832 => std_logic_vector(to_unsigned(2, 8)),
			6833 => std_logic_vector(to_unsigned(4, 8)),
			6834 => std_logic_vector(to_unsigned(181, 8)),
			6835 => std_logic_vector(to_unsigned(10, 8)),
			6836 => std_logic_vector(to_unsigned(255, 8)),
			6837 => std_logic_vector(to_unsigned(123, 8)),
			6838 => std_logic_vector(to_unsigned(153, 8)),
			6839 => std_logic_vector(to_unsigned(91, 8)),
			6840 => std_logic_vector(to_unsigned(65, 8)),
			6841 => std_logic_vector(to_unsigned(23, 8)),
			6842 => std_logic_vector(to_unsigned(159, 8)),
			6843 => std_logic_vector(to_unsigned(26, 8)),
			6844 => std_logic_vector(to_unsigned(71, 8)),
			6845 => std_logic_vector(to_unsigned(7, 8)),
			6846 => std_logic_vector(to_unsigned(88, 8)),
			6847 => std_logic_vector(to_unsigned(131, 8)),
			6848 => std_logic_vector(to_unsigned(79, 8)),
			6849 => std_logic_vector(to_unsigned(233, 8)),
			6850 => std_logic_vector(to_unsigned(54, 8)),
			6851 => std_logic_vector(to_unsigned(244, 8)),
			6852 => std_logic_vector(to_unsigned(207, 8)),
			6853 => std_logic_vector(to_unsigned(43, 8)),
			6854 => std_logic_vector(to_unsigned(68, 8)),
			6855 => std_logic_vector(to_unsigned(246, 8)),
			6856 => std_logic_vector(to_unsigned(241, 8)),
			6857 => std_logic_vector(to_unsigned(134, 8)),
			6858 => std_logic_vector(to_unsigned(237, 8)),
			6859 => std_logic_vector(to_unsigned(36, 8)),
			6860 => std_logic_vector(to_unsigned(101, 8)),
			6861 => std_logic_vector(to_unsigned(157, 8)),
			6862 => std_logic_vector(to_unsigned(233, 8)),
			6863 => std_logic_vector(to_unsigned(56, 8)),
			6864 => std_logic_vector(to_unsigned(117, 8)),
			6865 => std_logic_vector(to_unsigned(192, 8)),
			6866 => std_logic_vector(to_unsigned(173, 8)),
			6867 => std_logic_vector(to_unsigned(156, 8)),
			6868 => std_logic_vector(to_unsigned(189, 8)),
			6869 => std_logic_vector(to_unsigned(31, 8)),
			6870 => std_logic_vector(to_unsigned(94, 8)),
			6871 => std_logic_vector(to_unsigned(45, 8)),
			6872 => std_logic_vector(to_unsigned(186, 8)),
			6873 => std_logic_vector(to_unsigned(215, 8)),
			6874 => std_logic_vector(to_unsigned(131, 8)),
			6875 => std_logic_vector(to_unsigned(152, 8)),
			6876 => std_logic_vector(to_unsigned(243, 8)),
			6877 => std_logic_vector(to_unsigned(253, 8)),
			6878 => std_logic_vector(to_unsigned(242, 8)),
			6879 => std_logic_vector(to_unsigned(185, 8)),
			6880 => std_logic_vector(to_unsigned(201, 8)),
			6881 => std_logic_vector(to_unsigned(218, 8)),
			6882 => std_logic_vector(to_unsigned(103, 8)),
			6883 => std_logic_vector(to_unsigned(228, 8)),
			6884 => std_logic_vector(to_unsigned(155, 8)),
			6885 => std_logic_vector(to_unsigned(26, 8)),
			6886 => std_logic_vector(to_unsigned(160, 8)),
			6887 => std_logic_vector(to_unsigned(108, 8)),
			6888 => std_logic_vector(to_unsigned(36, 8)),
			6889 => std_logic_vector(to_unsigned(132, 8)),
			6890 => std_logic_vector(to_unsigned(117, 8)),
			6891 => std_logic_vector(to_unsigned(13, 8)),
			6892 => std_logic_vector(to_unsigned(218, 8)),
			6893 => std_logic_vector(to_unsigned(168, 8)),
			6894 => std_logic_vector(to_unsigned(176, 8)),
			6895 => std_logic_vector(to_unsigned(6, 8)),
			6896 => std_logic_vector(to_unsigned(45, 8)),
			6897 => std_logic_vector(to_unsigned(196, 8)),
			6898 => std_logic_vector(to_unsigned(228, 8)),
			6899 => std_logic_vector(to_unsigned(145, 8)),
			6900 => std_logic_vector(to_unsigned(21, 8)),
			6901 => std_logic_vector(to_unsigned(196, 8)),
			6902 => std_logic_vector(to_unsigned(240, 8)),
			6903 => std_logic_vector(to_unsigned(84, 8)),
			6904 => std_logic_vector(to_unsigned(26, 8)),
			6905 => std_logic_vector(to_unsigned(118, 8)),
			6906 => std_logic_vector(to_unsigned(138, 8)),
			6907 => std_logic_vector(to_unsigned(7, 8)),
			6908 => std_logic_vector(to_unsigned(77, 8)),
			6909 => std_logic_vector(to_unsigned(14, 8)),
			6910 => std_logic_vector(to_unsigned(62, 8)),
			6911 => std_logic_vector(to_unsigned(63, 8)),
			6912 => std_logic_vector(to_unsigned(87, 8)),
			6913 => std_logic_vector(to_unsigned(72, 8)),
			6914 => std_logic_vector(to_unsigned(138, 8)),
			6915 => std_logic_vector(to_unsigned(191, 8)),
			6916 => std_logic_vector(to_unsigned(179, 8)),
			6917 => std_logic_vector(to_unsigned(8, 8)),
			6918 => std_logic_vector(to_unsigned(222, 8)),
			6919 => std_logic_vector(to_unsigned(123, 8)),
			6920 => std_logic_vector(to_unsigned(93, 8)),
			6921 => std_logic_vector(to_unsigned(11, 8)),
			6922 => std_logic_vector(to_unsigned(142, 8)),
			6923 => std_logic_vector(to_unsigned(222, 8)),
			6924 => std_logic_vector(to_unsigned(56, 8)),
			6925 => std_logic_vector(to_unsigned(115, 8)),
			6926 => std_logic_vector(to_unsigned(27, 8)),
			6927 => std_logic_vector(to_unsigned(193, 8)),
			6928 => std_logic_vector(to_unsigned(233, 8)),
			6929 => std_logic_vector(to_unsigned(112, 8)),
			6930 => std_logic_vector(to_unsigned(63, 8)),
			6931 => std_logic_vector(to_unsigned(226, 8)),
			6932 => std_logic_vector(to_unsigned(200, 8)),
			6933 => std_logic_vector(to_unsigned(220, 8)),
			6934 => std_logic_vector(to_unsigned(208, 8)),
			6935 => std_logic_vector(to_unsigned(12, 8)),
			6936 => std_logic_vector(to_unsigned(126, 8)),
			6937 => std_logic_vector(to_unsigned(242, 8)),
			6938 => std_logic_vector(to_unsigned(163, 8)),
			6939 => std_logic_vector(to_unsigned(13, 8)),
			6940 => std_logic_vector(to_unsigned(194, 8)),
			6941 => std_logic_vector(to_unsigned(16, 8)),
			6942 => std_logic_vector(to_unsigned(208, 8)),
			6943 => std_logic_vector(to_unsigned(189, 8)),
			6944 => std_logic_vector(to_unsigned(148, 8)),
			6945 => std_logic_vector(to_unsigned(18, 8)),
			6946 => std_logic_vector(to_unsigned(144, 8)),
			6947 => std_logic_vector(to_unsigned(161, 8)),
			6948 => std_logic_vector(to_unsigned(212, 8)),
			6949 => std_logic_vector(to_unsigned(147, 8)),
			6950 => std_logic_vector(to_unsigned(65, 8)),
			6951 => std_logic_vector(to_unsigned(7, 8)),
			6952 => std_logic_vector(to_unsigned(173, 8)),
			6953 => std_logic_vector(to_unsigned(165, 8)),
			6954 => std_logic_vector(to_unsigned(129, 8)),
			6955 => std_logic_vector(to_unsigned(109, 8)),
			6956 => std_logic_vector(to_unsigned(71, 8)),
			6957 => std_logic_vector(to_unsigned(170, 8)),
			6958 => std_logic_vector(to_unsigned(159, 8)),
			6959 => std_logic_vector(to_unsigned(134, 8)),
			6960 => std_logic_vector(to_unsigned(160, 8)),
			6961 => std_logic_vector(to_unsigned(239, 8)),
			6962 => std_logic_vector(to_unsigned(216, 8)),
			6963 => std_logic_vector(to_unsigned(236, 8)),
			6964 => std_logic_vector(to_unsigned(141, 8)),
			6965 => std_logic_vector(to_unsigned(191, 8)),
			6966 => std_logic_vector(to_unsigned(154, 8)),
			6967 => std_logic_vector(to_unsigned(174, 8)),
			6968 => std_logic_vector(to_unsigned(199, 8)),
			6969 => std_logic_vector(to_unsigned(236, 8)),
			6970 => std_logic_vector(to_unsigned(136, 8)),
			6971 => std_logic_vector(to_unsigned(236, 8)),
			6972 => std_logic_vector(to_unsigned(132, 8)),
			6973 => std_logic_vector(to_unsigned(32, 8)),
			6974 => std_logic_vector(to_unsigned(101, 8)),
			6975 => std_logic_vector(to_unsigned(118, 8)),
			6976 => std_logic_vector(to_unsigned(43, 8)),
			6977 => std_logic_vector(to_unsigned(217, 8)),
			6978 => std_logic_vector(to_unsigned(235, 8)),
			6979 => std_logic_vector(to_unsigned(152, 8)),
			6980 => std_logic_vector(to_unsigned(102, 8)),
			6981 => std_logic_vector(to_unsigned(213, 8)),
			6982 => std_logic_vector(to_unsigned(42, 8)),
			6983 => std_logic_vector(to_unsigned(176, 8)),
			6984 => std_logic_vector(to_unsigned(3, 8)),
			6985 => std_logic_vector(to_unsigned(133, 8)),
			6986 => std_logic_vector(to_unsigned(232, 8)),
			6987 => std_logic_vector(to_unsigned(249, 8)),
			6988 => std_logic_vector(to_unsigned(85, 8)),
			6989 => std_logic_vector(to_unsigned(187, 8)),
			6990 => std_logic_vector(to_unsigned(206, 8)),
			6991 => std_logic_vector(to_unsigned(49, 8)),
			6992 => std_logic_vector(to_unsigned(170, 8)),
			6993 => std_logic_vector(to_unsigned(58, 8)),
			6994 => std_logic_vector(to_unsigned(10, 8)),
			6995 => std_logic_vector(to_unsigned(185, 8)),
			6996 => std_logic_vector(to_unsigned(94, 8)),
			6997 => std_logic_vector(to_unsigned(189, 8)),
			6998 => std_logic_vector(to_unsigned(134, 8)),
			6999 => std_logic_vector(to_unsigned(198, 8)),
			7000 => std_logic_vector(to_unsigned(188, 8)),
			7001 => std_logic_vector(to_unsigned(13, 8)),
			7002 => std_logic_vector(to_unsigned(136, 8)),
			7003 => std_logic_vector(to_unsigned(67, 8)),
			7004 => std_logic_vector(to_unsigned(189, 8)),
			7005 => std_logic_vector(to_unsigned(118, 8)),
			7006 => std_logic_vector(to_unsigned(59, 8)),
			7007 => std_logic_vector(to_unsigned(63, 8)),
			7008 => std_logic_vector(to_unsigned(83, 8)),
			7009 => std_logic_vector(to_unsigned(98, 8)),
			7010 => std_logic_vector(to_unsigned(230, 8)),
			7011 => std_logic_vector(to_unsigned(5, 8)),
			7012 => std_logic_vector(to_unsigned(179, 8)),
			7013 => std_logic_vector(to_unsigned(187, 8)),
			7014 => std_logic_vector(to_unsigned(65, 8)),
			7015 => std_logic_vector(to_unsigned(7, 8)),
			7016 => std_logic_vector(to_unsigned(30, 8)),
			7017 => std_logic_vector(to_unsigned(10, 8)),
			7018 => std_logic_vector(to_unsigned(73, 8)),
			7019 => std_logic_vector(to_unsigned(98, 8)),
			7020 => std_logic_vector(to_unsigned(254, 8)),
			7021 => std_logic_vector(to_unsigned(251, 8)),
			7022 => std_logic_vector(to_unsigned(95, 8)),
			7023 => std_logic_vector(to_unsigned(154, 8)),
			7024 => std_logic_vector(to_unsigned(20, 8)),
			7025 => std_logic_vector(to_unsigned(174, 8)),
			7026 => std_logic_vector(to_unsigned(175, 8)),
			7027 => std_logic_vector(to_unsigned(132, 8)),
			7028 => std_logic_vector(to_unsigned(139, 8)),
			7029 => std_logic_vector(to_unsigned(85, 8)),
			7030 => std_logic_vector(to_unsigned(93, 8)),
			7031 => std_logic_vector(to_unsigned(159, 8)),
			7032 => std_logic_vector(to_unsigned(188, 8)),
			7033 => std_logic_vector(to_unsigned(251, 8)),
			7034 => std_logic_vector(to_unsigned(16, 8)),
			7035 => std_logic_vector(to_unsigned(238, 8)),
			7036 => std_logic_vector(to_unsigned(218, 8)),
			7037 => std_logic_vector(to_unsigned(10, 8)),
			7038 => std_logic_vector(to_unsigned(255, 8)),
			7039 => std_logic_vector(to_unsigned(216, 8)),
			7040 => std_logic_vector(to_unsigned(127, 8)),
			7041 => std_logic_vector(to_unsigned(84, 8)),
			7042 => std_logic_vector(to_unsigned(89, 8)),
			7043 => std_logic_vector(to_unsigned(98, 8)),
			7044 => std_logic_vector(to_unsigned(212, 8)),
			7045 => std_logic_vector(to_unsigned(48, 8)),
			7046 => std_logic_vector(to_unsigned(239, 8)),
			7047 => std_logic_vector(to_unsigned(235, 8)),
			7048 => std_logic_vector(to_unsigned(219, 8)),
			7049 => std_logic_vector(to_unsigned(99, 8)),
			7050 => std_logic_vector(to_unsigned(234, 8)),
			7051 => std_logic_vector(to_unsigned(204, 8)),
			7052 => std_logic_vector(to_unsigned(194, 8)),
			7053 => std_logic_vector(to_unsigned(40, 8)),
			7054 => std_logic_vector(to_unsigned(76, 8)),
			7055 => std_logic_vector(to_unsigned(246, 8)),
			7056 => std_logic_vector(to_unsigned(238, 8)),
			7057 => std_logic_vector(to_unsigned(48, 8)),
			7058 => std_logic_vector(to_unsigned(184, 8)),
			7059 => std_logic_vector(to_unsigned(214, 8)),
			7060 => std_logic_vector(to_unsigned(37, 8)),
			7061 => std_logic_vector(to_unsigned(42, 8)),
			7062 => std_logic_vector(to_unsigned(27, 8)),
			7063 => std_logic_vector(to_unsigned(82, 8)),
			7064 => std_logic_vector(to_unsigned(211, 8)),
			7065 => std_logic_vector(to_unsigned(83, 8)),
			7066 => std_logic_vector(to_unsigned(33, 8)),
			7067 => std_logic_vector(to_unsigned(189, 8)),
			7068 => std_logic_vector(to_unsigned(122, 8)),
			7069 => std_logic_vector(to_unsigned(242, 8)),
			7070 => std_logic_vector(to_unsigned(31, 8)),
			7071 => std_logic_vector(to_unsigned(233, 8)),
			7072 => std_logic_vector(to_unsigned(40, 8)),
			7073 => std_logic_vector(to_unsigned(159, 8)),
			7074 => std_logic_vector(to_unsigned(82, 8)),
			7075 => std_logic_vector(to_unsigned(42, 8)),
			7076 => std_logic_vector(to_unsigned(60, 8)),
			7077 => std_logic_vector(to_unsigned(189, 8)),
			7078 => std_logic_vector(to_unsigned(228, 8)),
			7079 => std_logic_vector(to_unsigned(2, 8)),
			7080 => std_logic_vector(to_unsigned(251, 8)),
			7081 => std_logic_vector(to_unsigned(179, 8)),
			7082 => std_logic_vector(to_unsigned(116, 8)),
			7083 => std_logic_vector(to_unsigned(245, 8)),
			7084 => std_logic_vector(to_unsigned(220, 8)),
			7085 => std_logic_vector(to_unsigned(118, 8)),
			7086 => std_logic_vector(to_unsigned(205, 8)),
			7087 => std_logic_vector(to_unsigned(75, 8)),
			7088 => std_logic_vector(to_unsigned(186, 8)),
			7089 => std_logic_vector(to_unsigned(93, 8)),
			7090 => std_logic_vector(to_unsigned(57, 8)),
			7091 => std_logic_vector(to_unsigned(145, 8)),
			7092 => std_logic_vector(to_unsigned(215, 8)),
			7093 => std_logic_vector(to_unsigned(81, 8)),
			7094 => std_logic_vector(to_unsigned(225, 8)),
			7095 => std_logic_vector(to_unsigned(236, 8)),
			7096 => std_logic_vector(to_unsigned(200, 8)),
			7097 => std_logic_vector(to_unsigned(42, 8)),
			7098 => std_logic_vector(to_unsigned(116, 8)),
			7099 => std_logic_vector(to_unsigned(97, 8)),
			7100 => std_logic_vector(to_unsigned(244, 8)),
			7101 => std_logic_vector(to_unsigned(243, 8)),
			7102 => std_logic_vector(to_unsigned(140, 8)),
			7103 => std_logic_vector(to_unsigned(77, 8)),
			7104 => std_logic_vector(to_unsigned(60, 8)),
			7105 => std_logic_vector(to_unsigned(204, 8)),
			7106 => std_logic_vector(to_unsigned(166, 8)),
			7107 => std_logic_vector(to_unsigned(151, 8)),
			7108 => std_logic_vector(to_unsigned(231, 8)),
			7109 => std_logic_vector(to_unsigned(254, 8)),
			7110 => std_logic_vector(to_unsigned(174, 8)),
			7111 => std_logic_vector(to_unsigned(160, 8)),
			7112 => std_logic_vector(to_unsigned(62, 8)),
			7113 => std_logic_vector(to_unsigned(128, 8)),
			7114 => std_logic_vector(to_unsigned(199, 8)),
			7115 => std_logic_vector(to_unsigned(141, 8)),
			7116 => std_logic_vector(to_unsigned(224, 8)),
			7117 => std_logic_vector(to_unsigned(244, 8)),
			7118 => std_logic_vector(to_unsigned(42, 8)),
			7119 => std_logic_vector(to_unsigned(230, 8)),
			7120 => std_logic_vector(to_unsigned(65, 8)),
			7121 => std_logic_vector(to_unsigned(187, 8)),
			7122 => std_logic_vector(to_unsigned(244, 8)),
			7123 => std_logic_vector(to_unsigned(72, 8)),
			7124 => std_logic_vector(to_unsigned(63, 8)),
			7125 => std_logic_vector(to_unsigned(87, 8)),
			7126 => std_logic_vector(to_unsigned(249, 8)),
			7127 => std_logic_vector(to_unsigned(160, 8)),
			7128 => std_logic_vector(to_unsigned(137, 8)),
			7129 => std_logic_vector(to_unsigned(151, 8)),
			7130 => std_logic_vector(to_unsigned(185, 8)),
			7131 => std_logic_vector(to_unsigned(82, 8)),
			7132 => std_logic_vector(to_unsigned(51, 8)),
			7133 => std_logic_vector(to_unsigned(83, 8)),
			7134 => std_logic_vector(to_unsigned(135, 8)),
			7135 => std_logic_vector(to_unsigned(34, 8)),
			7136 => std_logic_vector(to_unsigned(220, 8)),
			7137 => std_logic_vector(to_unsigned(138, 8)),
			7138 => std_logic_vector(to_unsigned(138, 8)),
			7139 => std_logic_vector(to_unsigned(180, 8)),
			7140 => std_logic_vector(to_unsigned(159, 8)),
			7141 => std_logic_vector(to_unsigned(10, 8)),
			7142 => std_logic_vector(to_unsigned(219, 8)),
			7143 => std_logic_vector(to_unsigned(53, 8)),
			7144 => std_logic_vector(to_unsigned(196, 8)),
			7145 => std_logic_vector(to_unsigned(249, 8)),
			7146 => std_logic_vector(to_unsigned(60, 8)),
			7147 => std_logic_vector(to_unsigned(33, 8)),
			7148 => std_logic_vector(to_unsigned(143, 8)),
			7149 => std_logic_vector(to_unsigned(228, 8)),
			7150 => std_logic_vector(to_unsigned(228, 8)),
			7151 => std_logic_vector(to_unsigned(142, 8)),
			7152 => std_logic_vector(to_unsigned(236, 8)),
			7153 => std_logic_vector(to_unsigned(172, 8)),
			7154 => std_logic_vector(to_unsigned(133, 8)),
			7155 => std_logic_vector(to_unsigned(117, 8)),
			7156 => std_logic_vector(to_unsigned(183, 8)),
			7157 => std_logic_vector(to_unsigned(162, 8)),
			7158 => std_logic_vector(to_unsigned(60, 8)),
			7159 => std_logic_vector(to_unsigned(227, 8)),
			7160 => std_logic_vector(to_unsigned(254, 8)),
			7161 => std_logic_vector(to_unsigned(245, 8)),
			7162 => std_logic_vector(to_unsigned(50, 8)),
			7163 => std_logic_vector(to_unsigned(142, 8)),
			7164 => std_logic_vector(to_unsigned(61, 8)),
			7165 => std_logic_vector(to_unsigned(28, 8)),
			7166 => std_logic_vector(to_unsigned(86, 8)),
			7167 => std_logic_vector(to_unsigned(137, 8)),
			7168 => std_logic_vector(to_unsigned(152, 8)),
			7169 => std_logic_vector(to_unsigned(235, 8)),
			7170 => std_logic_vector(to_unsigned(213, 8)),
			7171 => std_logic_vector(to_unsigned(137, 8)),
			7172 => std_logic_vector(to_unsigned(220, 8)),
			7173 => std_logic_vector(to_unsigned(231, 8)),
			7174 => std_logic_vector(to_unsigned(173, 8)),
			7175 => std_logic_vector(to_unsigned(220, 8)),
			7176 => std_logic_vector(to_unsigned(197, 8)),
			7177 => std_logic_vector(to_unsigned(247, 8)),
			7178 => std_logic_vector(to_unsigned(142, 8)),
			7179 => std_logic_vector(to_unsigned(208, 8)),
			7180 => std_logic_vector(to_unsigned(120, 8)),
			7181 => std_logic_vector(to_unsigned(177, 8)),
			7182 => std_logic_vector(to_unsigned(178, 8)),
			7183 => std_logic_vector(to_unsigned(2, 8)),
			7184 => std_logic_vector(to_unsigned(175, 8)),
			7185 => std_logic_vector(to_unsigned(171, 8)),
			7186 => std_logic_vector(to_unsigned(164, 8)),
			7187 => std_logic_vector(to_unsigned(65, 8)),
			7188 => std_logic_vector(to_unsigned(115, 8)),
			7189 => std_logic_vector(to_unsigned(27, 8)),
			7190 => std_logic_vector(to_unsigned(185, 8)),
			7191 => std_logic_vector(to_unsigned(134, 8)),
			7192 => std_logic_vector(to_unsigned(236, 8)),
			7193 => std_logic_vector(to_unsigned(167, 8)),
			7194 => std_logic_vector(to_unsigned(225, 8)),
			7195 => std_logic_vector(to_unsigned(120, 8)),
			7196 => std_logic_vector(to_unsigned(102, 8)),
			7197 => std_logic_vector(to_unsigned(186, 8)),
			7198 => std_logic_vector(to_unsigned(157, 8)),
			7199 => std_logic_vector(to_unsigned(159, 8)),
			7200 => std_logic_vector(to_unsigned(242, 8)),
			7201 => std_logic_vector(to_unsigned(14, 8)),
			7202 => std_logic_vector(to_unsigned(153, 8)),
			7203 => std_logic_vector(to_unsigned(193, 8)),
			7204 => std_logic_vector(to_unsigned(161, 8)),
			7205 => std_logic_vector(to_unsigned(248, 8)),
			7206 => std_logic_vector(to_unsigned(11, 8)),
			7207 => std_logic_vector(to_unsigned(134, 8)),
			7208 => std_logic_vector(to_unsigned(125, 8)),
			7209 => std_logic_vector(to_unsigned(198, 8)),
			7210 => std_logic_vector(to_unsigned(211, 8)),
			7211 => std_logic_vector(to_unsigned(54, 8)),
			7212 => std_logic_vector(to_unsigned(146, 8)),
			7213 => std_logic_vector(to_unsigned(147, 8)),
			7214 => std_logic_vector(to_unsigned(154, 8)),
			7215 => std_logic_vector(to_unsigned(79, 8)),
			7216 => std_logic_vector(to_unsigned(45, 8)),
			7217 => std_logic_vector(to_unsigned(118, 8)),
			7218 => std_logic_vector(to_unsigned(186, 8)),
			7219 => std_logic_vector(to_unsigned(5, 8)),
			7220 => std_logic_vector(to_unsigned(227, 8)),
			7221 => std_logic_vector(to_unsigned(12, 8)),
			7222 => std_logic_vector(to_unsigned(43, 8)),
			7223 => std_logic_vector(to_unsigned(38, 8)),
			7224 => std_logic_vector(to_unsigned(60, 8)),
			7225 => std_logic_vector(to_unsigned(14, 8)),
			7226 => std_logic_vector(to_unsigned(162, 8)),
			7227 => std_logic_vector(to_unsigned(117, 8)),
			7228 => std_logic_vector(to_unsigned(219, 8)),
			7229 => std_logic_vector(to_unsigned(9, 8)),
			7230 => std_logic_vector(to_unsigned(173, 8)),
			7231 => std_logic_vector(to_unsigned(172, 8)),
			7232 => std_logic_vector(to_unsigned(120, 8)),
			7233 => std_logic_vector(to_unsigned(14, 8)),
			7234 => std_logic_vector(to_unsigned(157, 8)),
			7235 => std_logic_vector(to_unsigned(73, 8)),
			7236 => std_logic_vector(to_unsigned(219, 8)),
			7237 => std_logic_vector(to_unsigned(23, 8)),
			7238 => std_logic_vector(to_unsigned(38, 8)),
			7239 => std_logic_vector(to_unsigned(184, 8)),
			7240 => std_logic_vector(to_unsigned(206, 8)),
			7241 => std_logic_vector(to_unsigned(70, 8)),
			7242 => std_logic_vector(to_unsigned(248, 8)),
			7243 => std_logic_vector(to_unsigned(84, 8)),
			7244 => std_logic_vector(to_unsigned(16, 8)),
			7245 => std_logic_vector(to_unsigned(248, 8)),
			7246 => std_logic_vector(to_unsigned(239, 8)),
			7247 => std_logic_vector(to_unsigned(12, 8)),
			7248 => std_logic_vector(to_unsigned(75, 8)),
			7249 => std_logic_vector(to_unsigned(8, 8)),
			7250 => std_logic_vector(to_unsigned(180, 8)),
			7251 => std_logic_vector(to_unsigned(68, 8)),
			7252 => std_logic_vector(to_unsigned(48, 8)),
			7253 => std_logic_vector(to_unsigned(231, 8)),
			7254 => std_logic_vector(to_unsigned(56, 8)),
			7255 => std_logic_vector(to_unsigned(153, 8)),
			7256 => std_logic_vector(to_unsigned(253, 8)),
			7257 => std_logic_vector(to_unsigned(144, 8)),
			7258 => std_logic_vector(to_unsigned(77, 8)),
			7259 => std_logic_vector(to_unsigned(200, 8)),
			7260 => std_logic_vector(to_unsigned(204, 8)),
			7261 => std_logic_vector(to_unsigned(185, 8)),
			7262 => std_logic_vector(to_unsigned(52, 8)),
			7263 => std_logic_vector(to_unsigned(235, 8)),
			7264 => std_logic_vector(to_unsigned(189, 8)),
			7265 => std_logic_vector(to_unsigned(228, 8)),
			7266 => std_logic_vector(to_unsigned(15, 8)),
			7267 => std_logic_vector(to_unsigned(100, 8)),
			7268 => std_logic_vector(to_unsigned(0, 8)),
			7269 => std_logic_vector(to_unsigned(1, 8)),
			7270 => std_logic_vector(to_unsigned(243, 8)),
			7271 => std_logic_vector(to_unsigned(185, 8)),
			7272 => std_logic_vector(to_unsigned(3, 8)),
			7273 => std_logic_vector(to_unsigned(75, 8)),
			7274 => std_logic_vector(to_unsigned(49, 8)),
			7275 => std_logic_vector(to_unsigned(213, 8)),
			7276 => std_logic_vector(to_unsigned(4, 8)),
			7277 => std_logic_vector(to_unsigned(20, 8)),
			7278 => std_logic_vector(to_unsigned(99, 8)),
			7279 => std_logic_vector(to_unsigned(232, 8)),
			7280 => std_logic_vector(to_unsigned(231, 8)),
			7281 => std_logic_vector(to_unsigned(39, 8)),
			7282 => std_logic_vector(to_unsigned(8, 8)),
			7283 => std_logic_vector(to_unsigned(18, 8)),
			7284 => std_logic_vector(to_unsigned(20, 8)),
			7285 => std_logic_vector(to_unsigned(158, 8)),
			7286 => std_logic_vector(to_unsigned(65, 8)),
			7287 => std_logic_vector(to_unsigned(28, 8)),
			7288 => std_logic_vector(to_unsigned(169, 8)),
			7289 => std_logic_vector(to_unsigned(21, 8)),
			7290 => std_logic_vector(to_unsigned(176, 8)),
			7291 => std_logic_vector(to_unsigned(41, 8)),
			7292 => std_logic_vector(to_unsigned(94, 8)),
			7293 => std_logic_vector(to_unsigned(137, 8)),
			7294 => std_logic_vector(to_unsigned(116, 8)),
			7295 => std_logic_vector(to_unsigned(254, 8)),
			7296 => std_logic_vector(to_unsigned(104, 8)),
			7297 => std_logic_vector(to_unsigned(21, 8)),
			7298 => std_logic_vector(to_unsigned(10, 8)),
			7299 => std_logic_vector(to_unsigned(14, 8)),
			7300 => std_logic_vector(to_unsigned(113, 8)),
			7301 => std_logic_vector(to_unsigned(87, 8)),
			7302 => std_logic_vector(to_unsigned(207, 8)),
			7303 => std_logic_vector(to_unsigned(122, 8)),
			7304 => std_logic_vector(to_unsigned(186, 8)),
			7305 => std_logic_vector(to_unsigned(244, 8)),
			7306 => std_logic_vector(to_unsigned(254, 8)),
			7307 => std_logic_vector(to_unsigned(120, 8)),
			7308 => std_logic_vector(to_unsigned(209, 8)),
			7309 => std_logic_vector(to_unsigned(53, 8)),
			7310 => std_logic_vector(to_unsigned(77, 8)),
			7311 => std_logic_vector(to_unsigned(235, 8)),
			7312 => std_logic_vector(to_unsigned(36, 8)),
			7313 => std_logic_vector(to_unsigned(109, 8)),
			7314 => std_logic_vector(to_unsigned(143, 8)),
			7315 => std_logic_vector(to_unsigned(91, 8)),
			7316 => std_logic_vector(to_unsigned(185, 8)),
			7317 => std_logic_vector(to_unsigned(59, 8)),
			7318 => std_logic_vector(to_unsigned(150, 8)),
			7319 => std_logic_vector(to_unsigned(172, 8)),
			7320 => std_logic_vector(to_unsigned(49, 8)),
			7321 => std_logic_vector(to_unsigned(13, 8)),
			7322 => std_logic_vector(to_unsigned(37, 8)),
			7323 => std_logic_vector(to_unsigned(71, 8)),
			7324 => std_logic_vector(to_unsigned(96, 8)),
			7325 => std_logic_vector(to_unsigned(103, 8)),
			7326 => std_logic_vector(to_unsigned(252, 8)),
			7327 => std_logic_vector(to_unsigned(237, 8)),
			7328 => std_logic_vector(to_unsigned(225, 8)),
			7329 => std_logic_vector(to_unsigned(117, 8)),
			7330 => std_logic_vector(to_unsigned(101, 8)),
			7331 => std_logic_vector(to_unsigned(7, 8)),
			7332 => std_logic_vector(to_unsigned(150, 8)),
			7333 => std_logic_vector(to_unsigned(184, 8)),
			7334 => std_logic_vector(to_unsigned(57, 8)),
			7335 => std_logic_vector(to_unsigned(250, 8)),
			7336 => std_logic_vector(to_unsigned(158, 8)),
			7337 => std_logic_vector(to_unsigned(20, 8)),
			7338 => std_logic_vector(to_unsigned(179, 8)),
			7339 => std_logic_vector(to_unsigned(201, 8)),
			7340 => std_logic_vector(to_unsigned(50, 8)),
			7341 => std_logic_vector(to_unsigned(36, 8)),
			7342 => std_logic_vector(to_unsigned(41, 8)),
			7343 => std_logic_vector(to_unsigned(253, 8)),
			7344 => std_logic_vector(to_unsigned(205, 8)),
			7345 => std_logic_vector(to_unsigned(4, 8)),
			7346 => std_logic_vector(to_unsigned(154, 8)),
			7347 => std_logic_vector(to_unsigned(40, 8)),
			7348 => std_logic_vector(to_unsigned(51, 8)),
			7349 => std_logic_vector(to_unsigned(188, 8)),
			7350 => std_logic_vector(to_unsigned(40, 8)),
			7351 => std_logic_vector(to_unsigned(227, 8)),
			7352 => std_logic_vector(to_unsigned(142, 8)),
			7353 => std_logic_vector(to_unsigned(147, 8)),
			7354 => std_logic_vector(to_unsigned(88, 8)),
			7355 => std_logic_vector(to_unsigned(146, 8)),
			7356 => std_logic_vector(to_unsigned(162, 8)),
			7357 => std_logic_vector(to_unsigned(101, 8)),
			7358 => std_logic_vector(to_unsigned(23, 8)),
			7359 => std_logic_vector(to_unsigned(81, 8)),
			7360 => std_logic_vector(to_unsigned(203, 8)),
			7361 => std_logic_vector(to_unsigned(182, 8)),
			7362 => std_logic_vector(to_unsigned(83, 8)),
			7363 => std_logic_vector(to_unsigned(69, 8)),
			7364 => std_logic_vector(to_unsigned(81, 8)),
			7365 => std_logic_vector(to_unsigned(192, 8)),
			7366 => std_logic_vector(to_unsigned(44, 8)),
			7367 => std_logic_vector(to_unsigned(77, 8)),
			7368 => std_logic_vector(to_unsigned(1, 8)),
			7369 => std_logic_vector(to_unsigned(198, 8)),
			7370 => std_logic_vector(to_unsigned(166, 8)),
			7371 => std_logic_vector(to_unsigned(149, 8)),
			7372 => std_logic_vector(to_unsigned(194, 8)),
			7373 => std_logic_vector(to_unsigned(198, 8)),
			7374 => std_logic_vector(to_unsigned(37, 8)),
			7375 => std_logic_vector(to_unsigned(25, 8)),
			7376 => std_logic_vector(to_unsigned(80, 8)),
			7377 => std_logic_vector(to_unsigned(214, 8)),
			7378 => std_logic_vector(to_unsigned(92, 8)),
			7379 => std_logic_vector(to_unsigned(168, 8)),
			7380 => std_logic_vector(to_unsigned(76, 8)),
			7381 => std_logic_vector(to_unsigned(255, 8)),
			7382 => std_logic_vector(to_unsigned(18, 8)),
			7383 => std_logic_vector(to_unsigned(250, 8)),
			7384 => std_logic_vector(to_unsigned(130, 8)),
			7385 => std_logic_vector(to_unsigned(249, 8)),
			7386 => std_logic_vector(to_unsigned(247, 8)),
			7387 => std_logic_vector(to_unsigned(254, 8)),
			7388 => std_logic_vector(to_unsigned(123, 8)),
			7389 => std_logic_vector(to_unsigned(53, 8)),
			7390 => std_logic_vector(to_unsigned(42, 8)),
			7391 => std_logic_vector(to_unsigned(100, 8)),
			7392 => std_logic_vector(to_unsigned(2, 8)),
			7393 => std_logic_vector(to_unsigned(210, 8)),
			7394 => std_logic_vector(to_unsigned(185, 8)),
			7395 => std_logic_vector(to_unsigned(245, 8)),
			7396 => std_logic_vector(to_unsigned(116, 8)),
			7397 => std_logic_vector(to_unsigned(168, 8)),
			7398 => std_logic_vector(to_unsigned(34, 8)),
			7399 => std_logic_vector(to_unsigned(188, 8)),
			7400 => std_logic_vector(to_unsigned(12, 8)),
			7401 => std_logic_vector(to_unsigned(122, 8)),
			7402 => std_logic_vector(to_unsigned(189, 8)),
			7403 => std_logic_vector(to_unsigned(15, 8)),
			7404 => std_logic_vector(to_unsigned(7, 8)),
			7405 => std_logic_vector(to_unsigned(61, 8)),
			7406 => std_logic_vector(to_unsigned(198, 8)),
			7407 => std_logic_vector(to_unsigned(37, 8)),
			7408 => std_logic_vector(to_unsigned(119, 8)),
			7409 => std_logic_vector(to_unsigned(35, 8)),
			7410 => std_logic_vector(to_unsigned(167, 8)),
			7411 => std_logic_vector(to_unsigned(210, 8)),
			7412 => std_logic_vector(to_unsigned(16, 8)),
			7413 => std_logic_vector(to_unsigned(8, 8)),
			7414 => std_logic_vector(to_unsigned(145, 8)),
			7415 => std_logic_vector(to_unsigned(105, 8)),
			7416 => std_logic_vector(to_unsigned(156, 8)),
			7417 => std_logic_vector(to_unsigned(209, 8)),
			7418 => std_logic_vector(to_unsigned(105, 8)),
			7419 => std_logic_vector(to_unsigned(70, 8)),
			7420 => std_logic_vector(to_unsigned(188, 8)),
			7421 => std_logic_vector(to_unsigned(228, 8)),
			7422 => std_logic_vector(to_unsigned(239, 8)),
			7423 => std_logic_vector(to_unsigned(134, 8)),
			7424 => std_logic_vector(to_unsigned(138, 8)),
			7425 => std_logic_vector(to_unsigned(167, 8)),
			7426 => std_logic_vector(to_unsigned(198, 8)),
			7427 => std_logic_vector(to_unsigned(88, 8)),
			7428 => std_logic_vector(to_unsigned(21, 8)),
			7429 => std_logic_vector(to_unsigned(144, 8)),
			7430 => std_logic_vector(to_unsigned(86, 8)),
			7431 => std_logic_vector(to_unsigned(31, 8)),
			7432 => std_logic_vector(to_unsigned(172, 8)),
			7433 => std_logic_vector(to_unsigned(160, 8)),
			7434 => std_logic_vector(to_unsigned(55, 8)),
			7435 => std_logic_vector(to_unsigned(160, 8)),
			7436 => std_logic_vector(to_unsigned(90, 8)),
			7437 => std_logic_vector(to_unsigned(136, 8)),
			7438 => std_logic_vector(to_unsigned(244, 8)),
			7439 => std_logic_vector(to_unsigned(28, 8)),
			7440 => std_logic_vector(to_unsigned(136, 8)),
			7441 => std_logic_vector(to_unsigned(209, 8)),
			7442 => std_logic_vector(to_unsigned(93, 8)),
			7443 => std_logic_vector(to_unsigned(31, 8)),
			7444 => std_logic_vector(to_unsigned(67, 8)),
			7445 => std_logic_vector(to_unsigned(252, 8)),
			7446 => std_logic_vector(to_unsigned(21, 8)),
			7447 => std_logic_vector(to_unsigned(44, 8)),
			7448 => std_logic_vector(to_unsigned(11, 8)),
			7449 => std_logic_vector(to_unsigned(55, 8)),
			7450 => std_logic_vector(to_unsigned(178, 8)),
			7451 => std_logic_vector(to_unsigned(156, 8)),
			7452 => std_logic_vector(to_unsigned(197, 8)),
			7453 => std_logic_vector(to_unsigned(210, 8)),
			7454 => std_logic_vector(to_unsigned(14, 8)),
			7455 => std_logic_vector(to_unsigned(57, 8)),
			7456 => std_logic_vector(to_unsigned(1, 8)),
			7457 => std_logic_vector(to_unsigned(210, 8)),
			7458 => std_logic_vector(to_unsigned(188, 8)),
			7459 => std_logic_vector(to_unsigned(132, 8)),
			7460 => std_logic_vector(to_unsigned(45, 8)),
			7461 => std_logic_vector(to_unsigned(94, 8)),
			7462 => std_logic_vector(to_unsigned(169, 8)),
			7463 => std_logic_vector(to_unsigned(249, 8)),
			7464 => std_logic_vector(to_unsigned(151, 8)),
			7465 => std_logic_vector(to_unsigned(22, 8)),
			7466 => std_logic_vector(to_unsigned(11, 8)),
			7467 => std_logic_vector(to_unsigned(110, 8)),
			7468 => std_logic_vector(to_unsigned(144, 8)),
			7469 => std_logic_vector(to_unsigned(212, 8)),
			7470 => std_logic_vector(to_unsigned(125, 8)),
			7471 => std_logic_vector(to_unsigned(150, 8)),
			7472 => std_logic_vector(to_unsigned(224, 8)),
			7473 => std_logic_vector(to_unsigned(228, 8)),
			7474 => std_logic_vector(to_unsigned(181, 8)),
			7475 => std_logic_vector(to_unsigned(195, 8)),
			7476 => std_logic_vector(to_unsigned(156, 8)),
			7477 => std_logic_vector(to_unsigned(149, 8)),
			7478 => std_logic_vector(to_unsigned(110, 8)),
			7479 => std_logic_vector(to_unsigned(101, 8)),
			7480 => std_logic_vector(to_unsigned(142, 8)),
			7481 => std_logic_vector(to_unsigned(101, 8)),
			7482 => std_logic_vector(to_unsigned(230, 8)),
			7483 => std_logic_vector(to_unsigned(213, 8)),
			7484 => std_logic_vector(to_unsigned(150, 8)),
			7485 => std_logic_vector(to_unsigned(240, 8)),
			7486 => std_logic_vector(to_unsigned(62, 8)),
			7487 => std_logic_vector(to_unsigned(238, 8)),
			7488 => std_logic_vector(to_unsigned(204, 8)),
			7489 => std_logic_vector(to_unsigned(110, 8)),
			7490 => std_logic_vector(to_unsigned(203, 8)),
			7491 => std_logic_vector(to_unsigned(221, 8)),
			7492 => std_logic_vector(to_unsigned(4, 8)),
			7493 => std_logic_vector(to_unsigned(97, 8)),
			7494 => std_logic_vector(to_unsigned(214, 8)),
			7495 => std_logic_vector(to_unsigned(3, 8)),
			7496 => std_logic_vector(to_unsigned(228, 8)),
			7497 => std_logic_vector(to_unsigned(109, 8)),
			7498 => std_logic_vector(to_unsigned(86, 8)),
			7499 => std_logic_vector(to_unsigned(110, 8)),
			7500 => std_logic_vector(to_unsigned(119, 8)),
			7501 => std_logic_vector(to_unsigned(15, 8)),
			7502 => std_logic_vector(to_unsigned(137, 8)),
			7503 => std_logic_vector(to_unsigned(27, 8)),
			7504 => std_logic_vector(to_unsigned(168, 8)),
			7505 => std_logic_vector(to_unsigned(95, 8)),
			7506 => std_logic_vector(to_unsigned(237, 8)),
			7507 => std_logic_vector(to_unsigned(17, 8)),
			7508 => std_logic_vector(to_unsigned(175, 8)),
			7509 => std_logic_vector(to_unsigned(123, 8)),
			7510 => std_logic_vector(to_unsigned(228, 8)),
			7511 => std_logic_vector(to_unsigned(81, 8)),
			7512 => std_logic_vector(to_unsigned(219, 8)),
			7513 => std_logic_vector(to_unsigned(90, 8)),
			7514 => std_logic_vector(to_unsigned(56, 8)),
			7515 => std_logic_vector(to_unsigned(84, 8)),
			7516 => std_logic_vector(to_unsigned(174, 8)),
			7517 => std_logic_vector(to_unsigned(231, 8)),
			7518 => std_logic_vector(to_unsigned(103, 8)),
			7519 => std_logic_vector(to_unsigned(205, 8)),
			7520 => std_logic_vector(to_unsigned(78, 8)),
			7521 => std_logic_vector(to_unsigned(71, 8)),
			7522 => std_logic_vector(to_unsigned(236, 8)),
			7523 => std_logic_vector(to_unsigned(123, 8)),
			7524 => std_logic_vector(to_unsigned(78, 8)),
			7525 => std_logic_vector(to_unsigned(217, 8)),
			7526 => std_logic_vector(to_unsigned(77, 8)),
			7527 => std_logic_vector(to_unsigned(156, 8)),
			7528 => std_logic_vector(to_unsigned(137, 8)),
			7529 => std_logic_vector(to_unsigned(97, 8)),
			7530 => std_logic_vector(to_unsigned(163, 8)),
			7531 => std_logic_vector(to_unsigned(6, 8)),
			7532 => std_logic_vector(to_unsigned(226, 8)),
			7533 => std_logic_vector(to_unsigned(187, 8)),
			7534 => std_logic_vector(to_unsigned(176, 8)),
			7535 => std_logic_vector(to_unsigned(233, 8)),
			7536 => std_logic_vector(to_unsigned(216, 8)),
			7537 => std_logic_vector(to_unsigned(20, 8)),
			7538 => std_logic_vector(to_unsigned(86, 8)),
			7539 => std_logic_vector(to_unsigned(70, 8)),
			7540 => std_logic_vector(to_unsigned(50, 8)),
			7541 => std_logic_vector(to_unsigned(39, 8)),
			7542 => std_logic_vector(to_unsigned(196, 8)),
			7543 => std_logic_vector(to_unsigned(58, 8)),
			7544 => std_logic_vector(to_unsigned(150, 8)),
			7545 => std_logic_vector(to_unsigned(194, 8)),
			7546 => std_logic_vector(to_unsigned(216, 8)),
			7547 => std_logic_vector(to_unsigned(159, 8)),
			7548 => std_logic_vector(to_unsigned(123, 8)),
			7549 => std_logic_vector(to_unsigned(67, 8)),
			7550 => std_logic_vector(to_unsigned(113, 8)),
			7551 => std_logic_vector(to_unsigned(78, 8)),
			7552 => std_logic_vector(to_unsigned(237, 8)),
			7553 => std_logic_vector(to_unsigned(100, 8)),
			7554 => std_logic_vector(to_unsigned(154, 8)),
			7555 => std_logic_vector(to_unsigned(12, 8)),
			7556 => std_logic_vector(to_unsigned(71, 8)),
			7557 => std_logic_vector(to_unsigned(156, 8)),
			7558 => std_logic_vector(to_unsigned(19, 8)),
			7559 => std_logic_vector(to_unsigned(197, 8)),
			7560 => std_logic_vector(to_unsigned(35, 8)),
			7561 => std_logic_vector(to_unsigned(5, 8)),
			7562 => std_logic_vector(to_unsigned(246, 8)),
			7563 => std_logic_vector(to_unsigned(247, 8)),
			7564 => std_logic_vector(to_unsigned(235, 8)),
			7565 => std_logic_vector(to_unsigned(143, 8)),
			7566 => std_logic_vector(to_unsigned(180, 8)),
			7567 => std_logic_vector(to_unsigned(209, 8)),
			7568 => std_logic_vector(to_unsigned(221, 8)),
			7569 => std_logic_vector(to_unsigned(192, 8)),
			7570 => std_logic_vector(to_unsigned(177, 8)),
			7571 => std_logic_vector(to_unsigned(197, 8)),
			7572 => std_logic_vector(to_unsigned(204, 8)),
			7573 => std_logic_vector(to_unsigned(254, 8)),
			7574 => std_logic_vector(to_unsigned(109, 8)),
			7575 => std_logic_vector(to_unsigned(130, 8)),
			7576 => std_logic_vector(to_unsigned(251, 8)),
			7577 => std_logic_vector(to_unsigned(187, 8)),
			7578 => std_logic_vector(to_unsigned(20, 8)),
			7579 => std_logic_vector(to_unsigned(89, 8)),
			7580 => std_logic_vector(to_unsigned(60, 8)),
			7581 => std_logic_vector(to_unsigned(220, 8)),
			7582 => std_logic_vector(to_unsigned(255, 8)),
			7583 => std_logic_vector(to_unsigned(25, 8)),
			7584 => std_logic_vector(to_unsigned(163, 8)),
			7585 => std_logic_vector(to_unsigned(203, 8)),
			7586 => std_logic_vector(to_unsigned(214, 8)),
			7587 => std_logic_vector(to_unsigned(192, 8)),
			7588 => std_logic_vector(to_unsigned(1, 8)),
			7589 => std_logic_vector(to_unsigned(227, 8)),
			7590 => std_logic_vector(to_unsigned(221, 8)),
			7591 => std_logic_vector(to_unsigned(107, 8)),
			7592 => std_logic_vector(to_unsigned(203, 8)),
			7593 => std_logic_vector(to_unsigned(19, 8)),
			7594 => std_logic_vector(to_unsigned(115, 8)),
			7595 => std_logic_vector(to_unsigned(119, 8)),
			7596 => std_logic_vector(to_unsigned(18, 8)),
			7597 => std_logic_vector(to_unsigned(77, 8)),
			7598 => std_logic_vector(to_unsigned(154, 8)),
			7599 => std_logic_vector(to_unsigned(120, 8)),
			7600 => std_logic_vector(to_unsigned(38, 8)),
			7601 => std_logic_vector(to_unsigned(122, 8)),
			7602 => std_logic_vector(to_unsigned(212, 8)),
			7603 => std_logic_vector(to_unsigned(223, 8)),
			7604 => std_logic_vector(to_unsigned(39, 8)),
			7605 => std_logic_vector(to_unsigned(72, 8)),
			7606 => std_logic_vector(to_unsigned(136, 8)),
			7607 => std_logic_vector(to_unsigned(142, 8)),
			7608 => std_logic_vector(to_unsigned(206, 8)),
			7609 => std_logic_vector(to_unsigned(130, 8)),
			7610 => std_logic_vector(to_unsigned(130, 8)),
			7611 => std_logic_vector(to_unsigned(120, 8)),
			7612 => std_logic_vector(to_unsigned(116, 8)),
			7613 => std_logic_vector(to_unsigned(155, 8)),
			7614 => std_logic_vector(to_unsigned(214, 8)),
			7615 => std_logic_vector(to_unsigned(255, 8)),
			7616 => std_logic_vector(to_unsigned(236, 8)),
			7617 => std_logic_vector(to_unsigned(61, 8)),
			7618 => std_logic_vector(to_unsigned(63, 8)),
			7619 => std_logic_vector(to_unsigned(162, 8)),
			7620 => std_logic_vector(to_unsigned(210, 8)),
			7621 => std_logic_vector(to_unsigned(75, 8)),
			7622 => std_logic_vector(to_unsigned(155, 8)),
			7623 => std_logic_vector(to_unsigned(42, 8)),
			7624 => std_logic_vector(to_unsigned(228, 8)),
			7625 => std_logic_vector(to_unsigned(187, 8)),
			7626 => std_logic_vector(to_unsigned(121, 8)),
			7627 => std_logic_vector(to_unsigned(201, 8)),
			7628 => std_logic_vector(to_unsigned(77, 8)),
			7629 => std_logic_vector(to_unsigned(102, 8)),
			7630 => std_logic_vector(to_unsigned(246, 8)),
			7631 => std_logic_vector(to_unsigned(17, 8)),
			7632 => std_logic_vector(to_unsigned(18, 8)),
			7633 => std_logic_vector(to_unsigned(43, 8)),
			7634 => std_logic_vector(to_unsigned(104, 8)),
			7635 => std_logic_vector(to_unsigned(51, 8)),
			7636 => std_logic_vector(to_unsigned(24, 8)),
			7637 => std_logic_vector(to_unsigned(120, 8)),
			7638 => std_logic_vector(to_unsigned(226, 8)),
			7639 => std_logic_vector(to_unsigned(196, 8)),
			7640 => std_logic_vector(to_unsigned(232, 8)),
			7641 => std_logic_vector(to_unsigned(145, 8)),
			7642 => std_logic_vector(to_unsigned(115, 8)),
			7643 => std_logic_vector(to_unsigned(39, 8)),
			7644 => std_logic_vector(to_unsigned(87, 8)),
			7645 => std_logic_vector(to_unsigned(210, 8)),
			7646 => std_logic_vector(to_unsigned(144, 8)),
			7647 => std_logic_vector(to_unsigned(151, 8)),
			7648 => std_logic_vector(to_unsigned(154, 8)),
			7649 => std_logic_vector(to_unsigned(77, 8)),
			7650 => std_logic_vector(to_unsigned(58, 8)),
			7651 => std_logic_vector(to_unsigned(234, 8)),
			7652 => std_logic_vector(to_unsigned(47, 8)),
			7653 => std_logic_vector(to_unsigned(193, 8)),
			7654 => std_logic_vector(to_unsigned(106, 8)),
			7655 => std_logic_vector(to_unsigned(25, 8)),
			7656 => std_logic_vector(to_unsigned(225, 8)),
			7657 => std_logic_vector(to_unsigned(231, 8)),
			7658 => std_logic_vector(to_unsigned(44, 8)),
			7659 => std_logic_vector(to_unsigned(137, 8)),
			7660 => std_logic_vector(to_unsigned(125, 8)),
			7661 => std_logic_vector(to_unsigned(115, 8)),
			7662 => std_logic_vector(to_unsigned(110, 8)),
			7663 => std_logic_vector(to_unsigned(156, 8)),
			7664 => std_logic_vector(to_unsigned(6, 8)),
			7665 => std_logic_vector(to_unsigned(226, 8)),
			7666 => std_logic_vector(to_unsigned(46, 8)),
			7667 => std_logic_vector(to_unsigned(68, 8)),
			7668 => std_logic_vector(to_unsigned(2, 8)),
			7669 => std_logic_vector(to_unsigned(27, 8)),
			7670 => std_logic_vector(to_unsigned(88, 8)),
			7671 => std_logic_vector(to_unsigned(176, 8)),
			7672 => std_logic_vector(to_unsigned(12, 8)),
			7673 => std_logic_vector(to_unsigned(40, 8)),
			7674 => std_logic_vector(to_unsigned(76, 8)),
			7675 => std_logic_vector(to_unsigned(220, 8)),
			7676 => std_logic_vector(to_unsigned(217, 8)),
			7677 => std_logic_vector(to_unsigned(183, 8)),
			7678 => std_logic_vector(to_unsigned(0, 8)),
			7679 => std_logic_vector(to_unsigned(116, 8)),
			7680 => std_logic_vector(to_unsigned(47, 8)),
			7681 => std_logic_vector(to_unsigned(105, 8)),
			7682 => std_logic_vector(to_unsigned(64, 8)),
			7683 => std_logic_vector(to_unsigned(176, 8)),
			7684 => std_logic_vector(to_unsigned(51, 8)),
			7685 => std_logic_vector(to_unsigned(34, 8)),
			7686 => std_logic_vector(to_unsigned(163, 8)),
			7687 => std_logic_vector(to_unsigned(62, 8)),
			7688 => std_logic_vector(to_unsigned(17, 8)),
			7689 => std_logic_vector(to_unsigned(206, 8)),
			7690 => std_logic_vector(to_unsigned(85, 8)),
			7691 => std_logic_vector(to_unsigned(82, 8)),
			7692 => std_logic_vector(to_unsigned(191, 8)),
			7693 => std_logic_vector(to_unsigned(231, 8)),
			7694 => std_logic_vector(to_unsigned(183, 8)),
			7695 => std_logic_vector(to_unsigned(142, 8)),
			7696 => std_logic_vector(to_unsigned(186, 8)),
			7697 => std_logic_vector(to_unsigned(26, 8)),
			7698 => std_logic_vector(to_unsigned(209, 8)),
			7699 => std_logic_vector(to_unsigned(253, 8)),
			7700 => std_logic_vector(to_unsigned(71, 8)),
			7701 => std_logic_vector(to_unsigned(145, 8)),
			7702 => std_logic_vector(to_unsigned(120, 8)),
			7703 => std_logic_vector(to_unsigned(228, 8)),
			7704 => std_logic_vector(to_unsigned(234, 8)),
			7705 => std_logic_vector(to_unsigned(47, 8)),
			7706 => std_logic_vector(to_unsigned(11, 8)),
			7707 => std_logic_vector(to_unsigned(86, 8)),
			7708 => std_logic_vector(to_unsigned(53, 8)),
			7709 => std_logic_vector(to_unsigned(75, 8)),
			7710 => std_logic_vector(to_unsigned(127, 8)),
			7711 => std_logic_vector(to_unsigned(196, 8)),
			7712 => std_logic_vector(to_unsigned(227, 8)),
			7713 => std_logic_vector(to_unsigned(237, 8)),
			7714 => std_logic_vector(to_unsigned(111, 8)),
			7715 => std_logic_vector(to_unsigned(168, 8)),
			7716 => std_logic_vector(to_unsigned(150, 8)),
			7717 => std_logic_vector(to_unsigned(126, 8)),
			7718 => std_logic_vector(to_unsigned(107, 8)),
			7719 => std_logic_vector(to_unsigned(155, 8)),
			7720 => std_logic_vector(to_unsigned(189, 8)),
			7721 => std_logic_vector(to_unsigned(96, 8)),
			7722 => std_logic_vector(to_unsigned(86, 8)),
			7723 => std_logic_vector(to_unsigned(106, 8)),
			7724 => std_logic_vector(to_unsigned(61, 8)),
			7725 => std_logic_vector(to_unsigned(118, 8)),
			7726 => std_logic_vector(to_unsigned(109, 8)),
			7727 => std_logic_vector(to_unsigned(122, 8)),
			7728 => std_logic_vector(to_unsigned(84, 8)),
			7729 => std_logic_vector(to_unsigned(75, 8)),
			7730 => std_logic_vector(to_unsigned(35, 8)),
			7731 => std_logic_vector(to_unsigned(77, 8)),
			7732 => std_logic_vector(to_unsigned(70, 8)),
			7733 => std_logic_vector(to_unsigned(49, 8)),
			7734 => std_logic_vector(to_unsigned(19, 8)),
			7735 => std_logic_vector(to_unsigned(233, 8)),
			7736 => std_logic_vector(to_unsigned(185, 8)),
			7737 => std_logic_vector(to_unsigned(157, 8)),
			7738 => std_logic_vector(to_unsigned(23, 8)),
			7739 => std_logic_vector(to_unsigned(55, 8)),
			7740 => std_logic_vector(to_unsigned(141, 8)),
			7741 => std_logic_vector(to_unsigned(150, 8)),
			7742 => std_logic_vector(to_unsigned(147, 8)),
			7743 => std_logic_vector(to_unsigned(126, 8)),
			7744 => std_logic_vector(to_unsigned(92, 8)),
			7745 => std_logic_vector(to_unsigned(9, 8)),
			7746 => std_logic_vector(to_unsigned(88, 8)),
			7747 => std_logic_vector(to_unsigned(113, 8)),
			7748 => std_logic_vector(to_unsigned(214, 8)),
			7749 => std_logic_vector(to_unsigned(132, 8)),
			7750 => std_logic_vector(to_unsigned(65, 8)),
			7751 => std_logic_vector(to_unsigned(92, 8)),
			7752 => std_logic_vector(to_unsigned(76, 8)),
			7753 => std_logic_vector(to_unsigned(23, 8)),
			7754 => std_logic_vector(to_unsigned(194, 8)),
			7755 => std_logic_vector(to_unsigned(170, 8)),
			7756 => std_logic_vector(to_unsigned(16, 8)),
			7757 => std_logic_vector(to_unsigned(53, 8)),
			7758 => std_logic_vector(to_unsigned(155, 8)),
			7759 => std_logic_vector(to_unsigned(217, 8)),
			7760 => std_logic_vector(to_unsigned(37, 8)),
			7761 => std_logic_vector(to_unsigned(230, 8)),
			7762 => std_logic_vector(to_unsigned(135, 8)),
			7763 => std_logic_vector(to_unsigned(143, 8)),
			7764 => std_logic_vector(to_unsigned(145, 8)),
			7765 => std_logic_vector(to_unsigned(92, 8)),
			7766 => std_logic_vector(to_unsigned(71, 8)),
			7767 => std_logic_vector(to_unsigned(252, 8)),
			7768 => std_logic_vector(to_unsigned(45, 8)),
			7769 => std_logic_vector(to_unsigned(133, 8)),
			7770 => std_logic_vector(to_unsigned(75, 8)),
			7771 => std_logic_vector(to_unsigned(180, 8)),
			7772 => std_logic_vector(to_unsigned(145, 8)),
			7773 => std_logic_vector(to_unsigned(222, 8)),
			7774 => std_logic_vector(to_unsigned(38, 8)),
			7775 => std_logic_vector(to_unsigned(140, 8)),
			7776 => std_logic_vector(to_unsigned(146, 8)),
			7777 => std_logic_vector(to_unsigned(190, 8)),
			7778 => std_logic_vector(to_unsigned(231, 8)),
			7779 => std_logic_vector(to_unsigned(125, 8)),
			7780 => std_logic_vector(to_unsigned(224, 8)),
			7781 => std_logic_vector(to_unsigned(236, 8)),
			7782 => std_logic_vector(to_unsigned(134, 8)),
			7783 => std_logic_vector(to_unsigned(189, 8)),
			7784 => std_logic_vector(to_unsigned(95, 8)),
			7785 => std_logic_vector(to_unsigned(213, 8)),
			7786 => std_logic_vector(to_unsigned(66, 8)),
			7787 => std_logic_vector(to_unsigned(7, 8)),
			7788 => std_logic_vector(to_unsigned(93, 8)),
			7789 => std_logic_vector(to_unsigned(143, 8)),
			7790 => std_logic_vector(to_unsigned(33, 8)),
			7791 => std_logic_vector(to_unsigned(254, 8)),
			7792 => std_logic_vector(to_unsigned(16, 8)),
			7793 => std_logic_vector(to_unsigned(206, 8)),
			7794 => std_logic_vector(to_unsigned(11, 8)),
			7795 => std_logic_vector(to_unsigned(162, 8)),
			7796 => std_logic_vector(to_unsigned(232, 8)),
			7797 => std_logic_vector(to_unsigned(159, 8)),
			7798 => std_logic_vector(to_unsigned(217, 8)),
			7799 => std_logic_vector(to_unsigned(102, 8)),
			7800 => std_logic_vector(to_unsigned(28, 8)),
			7801 => std_logic_vector(to_unsigned(180, 8)),
			7802 => std_logic_vector(to_unsigned(215, 8)),
			7803 => std_logic_vector(to_unsigned(25, 8)),
			7804 => std_logic_vector(to_unsigned(82, 8)),
			7805 => std_logic_vector(to_unsigned(197, 8)),
			7806 => std_logic_vector(to_unsigned(91, 8)),
			7807 => std_logic_vector(to_unsigned(239, 8)),
			7808 => std_logic_vector(to_unsigned(106, 8)),
			7809 => std_logic_vector(to_unsigned(239, 8)),
			7810 => std_logic_vector(to_unsigned(0, 8)),
			7811 => std_logic_vector(to_unsigned(129, 8)),
			7812 => std_logic_vector(to_unsigned(226, 8)),
			7813 => std_logic_vector(to_unsigned(245, 8)),
			7814 => std_logic_vector(to_unsigned(195, 8)),
			7815 => std_logic_vector(to_unsigned(62, 8)),
			7816 => std_logic_vector(to_unsigned(215, 8)),
			7817 => std_logic_vector(to_unsigned(87, 8)),
			7818 => std_logic_vector(to_unsigned(82, 8)),
			7819 => std_logic_vector(to_unsigned(178, 8)),
			7820 => std_logic_vector(to_unsigned(151, 8)),
			7821 => std_logic_vector(to_unsigned(104, 8)),
			7822 => std_logic_vector(to_unsigned(106, 8)),
			7823 => std_logic_vector(to_unsigned(53, 8)),
			7824 => std_logic_vector(to_unsigned(92, 8)),
			7825 => std_logic_vector(to_unsigned(17, 8)),
			7826 => std_logic_vector(to_unsigned(45, 8)),
			7827 => std_logic_vector(to_unsigned(101, 8)),
			7828 => std_logic_vector(to_unsigned(154, 8)),
			7829 => std_logic_vector(to_unsigned(240, 8)),
			7830 => std_logic_vector(to_unsigned(226, 8)),
			7831 => std_logic_vector(to_unsigned(114, 8)),
			7832 => std_logic_vector(to_unsigned(183, 8)),
			7833 => std_logic_vector(to_unsigned(126, 8)),
			7834 => std_logic_vector(to_unsigned(97, 8)),
			7835 => std_logic_vector(to_unsigned(243, 8)),
			7836 => std_logic_vector(to_unsigned(71, 8)),
			7837 => std_logic_vector(to_unsigned(113, 8)),
			7838 => std_logic_vector(to_unsigned(63, 8)),
			7839 => std_logic_vector(to_unsigned(60, 8)),
			7840 => std_logic_vector(to_unsigned(110, 8)),
			7841 => std_logic_vector(to_unsigned(80, 8)),
			7842 => std_logic_vector(to_unsigned(192, 8)),
			7843 => std_logic_vector(to_unsigned(135, 8)),
			7844 => std_logic_vector(to_unsigned(174, 8)),
			7845 => std_logic_vector(to_unsigned(59, 8)),
			7846 => std_logic_vector(to_unsigned(186, 8)),
			7847 => std_logic_vector(to_unsigned(217, 8)),
			7848 => std_logic_vector(to_unsigned(151, 8)),
			7849 => std_logic_vector(to_unsigned(189, 8)),
			7850 => std_logic_vector(to_unsigned(122, 8)),
			7851 => std_logic_vector(to_unsigned(47, 8)),
			7852 => std_logic_vector(to_unsigned(218, 8)),
			7853 => std_logic_vector(to_unsigned(123, 8)),
			7854 => std_logic_vector(to_unsigned(154, 8)),
			7855 => std_logic_vector(to_unsigned(159, 8)),
			7856 => std_logic_vector(to_unsigned(43, 8)),
			7857 => std_logic_vector(to_unsigned(183, 8)),
			7858 => std_logic_vector(to_unsigned(251, 8)),
			7859 => std_logic_vector(to_unsigned(252, 8)),
			7860 => std_logic_vector(to_unsigned(233, 8)),
			7861 => std_logic_vector(to_unsigned(220, 8)),
			7862 => std_logic_vector(to_unsigned(45, 8)),
			7863 => std_logic_vector(to_unsigned(156, 8)),
			7864 => std_logic_vector(to_unsigned(209, 8)),
			7865 => std_logic_vector(to_unsigned(10, 8)),
			7866 => std_logic_vector(to_unsigned(134, 8)),
			7867 => std_logic_vector(to_unsigned(149, 8)),
			7868 => std_logic_vector(to_unsigned(43, 8)),
			7869 => std_logic_vector(to_unsigned(35, 8)),
			7870 => std_logic_vector(to_unsigned(235, 8)),
			7871 => std_logic_vector(to_unsigned(246, 8)),
			7872 => std_logic_vector(to_unsigned(171, 8)),
			7873 => std_logic_vector(to_unsigned(243, 8)),
			7874 => std_logic_vector(to_unsigned(78, 8)),
			7875 => std_logic_vector(to_unsigned(197, 8)),
			7876 => std_logic_vector(to_unsigned(157, 8)),
			7877 => std_logic_vector(to_unsigned(197, 8)),
			7878 => std_logic_vector(to_unsigned(97, 8)),
			7879 => std_logic_vector(to_unsigned(102, 8)),
			7880 => std_logic_vector(to_unsigned(248, 8)),
			7881 => std_logic_vector(to_unsigned(76, 8)),
			7882 => std_logic_vector(to_unsigned(29, 8)),
			7883 => std_logic_vector(to_unsigned(130, 8)),
			7884 => std_logic_vector(to_unsigned(251, 8)),
			7885 => std_logic_vector(to_unsigned(222, 8)),
			7886 => std_logic_vector(to_unsigned(229, 8)),
			7887 => std_logic_vector(to_unsigned(22, 8)),
			7888 => std_logic_vector(to_unsigned(4, 8)),
			7889 => std_logic_vector(to_unsigned(166, 8)),
			7890 => std_logic_vector(to_unsigned(105, 8)),
			7891 => std_logic_vector(to_unsigned(83, 8)),
			7892 => std_logic_vector(to_unsigned(56, 8)),
			7893 => std_logic_vector(to_unsigned(161, 8)),
			7894 => std_logic_vector(to_unsigned(203, 8)),
			7895 => std_logic_vector(to_unsigned(63, 8)),
			7896 => std_logic_vector(to_unsigned(207, 8)),
			7897 => std_logic_vector(to_unsigned(247, 8)),
			7898 => std_logic_vector(to_unsigned(141, 8)),
			7899 => std_logic_vector(to_unsigned(45, 8)),
			7900 => std_logic_vector(to_unsigned(21, 8)),
			7901 => std_logic_vector(to_unsigned(141, 8)),
			7902 => std_logic_vector(to_unsigned(102, 8)),
			7903 => std_logic_vector(to_unsigned(196, 8)),
			7904 => std_logic_vector(to_unsigned(149, 8)),
			7905 => std_logic_vector(to_unsigned(118, 8)),
			7906 => std_logic_vector(to_unsigned(203, 8)),
			7907 => std_logic_vector(to_unsigned(100, 8)),
			7908 => std_logic_vector(to_unsigned(159, 8)),
			7909 => std_logic_vector(to_unsigned(243, 8)),
			7910 => std_logic_vector(to_unsigned(65, 8)),
			7911 => std_logic_vector(to_unsigned(42, 8)),
			7912 => std_logic_vector(to_unsigned(101, 8)),
			7913 => std_logic_vector(to_unsigned(191, 8)),
			7914 => std_logic_vector(to_unsigned(232, 8)),
			7915 => std_logic_vector(to_unsigned(98, 8)),
			7916 => std_logic_vector(to_unsigned(153, 8)),
			7917 => std_logic_vector(to_unsigned(127, 8)),
			7918 => std_logic_vector(to_unsigned(80, 8)),
			7919 => std_logic_vector(to_unsigned(255, 8)),
			7920 => std_logic_vector(to_unsigned(244, 8)),
			7921 => std_logic_vector(to_unsigned(138, 8)),
			7922 => std_logic_vector(to_unsigned(68, 8)),
			7923 => std_logic_vector(to_unsigned(32, 8)),
			7924 => std_logic_vector(to_unsigned(167, 8)),
			7925 => std_logic_vector(to_unsigned(50, 8)),
			7926 => std_logic_vector(to_unsigned(168, 8)),
			7927 => std_logic_vector(to_unsigned(165, 8)),
			7928 => std_logic_vector(to_unsigned(41, 8)),
			7929 => std_logic_vector(to_unsigned(37, 8)),
			7930 => std_logic_vector(to_unsigned(218, 8)),
			7931 => std_logic_vector(to_unsigned(212, 8)),
			7932 => std_logic_vector(to_unsigned(245, 8)),
			7933 => std_logic_vector(to_unsigned(76, 8)),
			7934 => std_logic_vector(to_unsigned(220, 8)),
			7935 => std_logic_vector(to_unsigned(9, 8)),
			7936 => std_logic_vector(to_unsigned(206, 8)),
			7937 => std_logic_vector(to_unsigned(94, 8)),
			7938 => std_logic_vector(to_unsigned(2, 8)),
			7939 => std_logic_vector(to_unsigned(30, 8)),
			7940 => std_logic_vector(to_unsigned(127, 8)),
			7941 => std_logic_vector(to_unsigned(77, 8)),
			7942 => std_logic_vector(to_unsigned(253, 8)),
			7943 => std_logic_vector(to_unsigned(190, 8)),
			7944 => std_logic_vector(to_unsigned(117, 8)),
			7945 => std_logic_vector(to_unsigned(1, 8)),
			7946 => std_logic_vector(to_unsigned(253, 8)),
			7947 => std_logic_vector(to_unsigned(157, 8)),
			7948 => std_logic_vector(to_unsigned(12, 8)),
			7949 => std_logic_vector(to_unsigned(217, 8)),
			7950 => std_logic_vector(to_unsigned(130, 8)),
			7951 => std_logic_vector(to_unsigned(107, 8)),
			7952 => std_logic_vector(to_unsigned(209, 8)),
			7953 => std_logic_vector(to_unsigned(130, 8)),
			7954 => std_logic_vector(to_unsigned(30, 8)),
			7955 => std_logic_vector(to_unsigned(148, 8)),
			7956 => std_logic_vector(to_unsigned(220, 8)),
			7957 => std_logic_vector(to_unsigned(16, 8)),
			7958 => std_logic_vector(to_unsigned(166, 8)),
			7959 => std_logic_vector(to_unsigned(71, 8)),
			7960 => std_logic_vector(to_unsigned(158, 8)),
			7961 => std_logic_vector(to_unsigned(107, 8)),
			7962 => std_logic_vector(to_unsigned(101, 8)),
			7963 => std_logic_vector(to_unsigned(218, 8)),
			7964 => std_logic_vector(to_unsigned(230, 8)),
			7965 => std_logic_vector(to_unsigned(54, 8)),
			7966 => std_logic_vector(to_unsigned(107, 8)),
			7967 => std_logic_vector(to_unsigned(6, 8)),
			7968 => std_logic_vector(to_unsigned(10, 8)),
			7969 => std_logic_vector(to_unsigned(244, 8)),
			7970 => std_logic_vector(to_unsigned(75, 8)),
			7971 => std_logic_vector(to_unsigned(189, 8)),
			7972 => std_logic_vector(to_unsigned(86, 8)),
			7973 => std_logic_vector(to_unsigned(123, 8)),
			7974 => std_logic_vector(to_unsigned(129, 8)),
			7975 => std_logic_vector(to_unsigned(95, 8)),
			7976 => std_logic_vector(to_unsigned(142, 8)),
			7977 => std_logic_vector(to_unsigned(3, 8)),
			7978 => std_logic_vector(to_unsigned(153, 8)),
			7979 => std_logic_vector(to_unsigned(97, 8)),
			7980 => std_logic_vector(to_unsigned(182, 8)),
			7981 => std_logic_vector(to_unsigned(138, 8)),
			7982 => std_logic_vector(to_unsigned(45, 8)),
			7983 => std_logic_vector(to_unsigned(12, 8)),
			7984 => std_logic_vector(to_unsigned(162, 8)),
			7985 => std_logic_vector(to_unsigned(155, 8)),
			7986 => std_logic_vector(to_unsigned(23, 8)),
			7987 => std_logic_vector(to_unsigned(167, 8)),
			7988 => std_logic_vector(to_unsigned(168, 8)),
			7989 => std_logic_vector(to_unsigned(161, 8)),
			7990 => std_logic_vector(to_unsigned(74, 8)),
			7991 => std_logic_vector(to_unsigned(57, 8)),
			7992 => std_logic_vector(to_unsigned(158, 8)),
			7993 => std_logic_vector(to_unsigned(158, 8)),
			7994 => std_logic_vector(to_unsigned(43, 8)),
			7995 => std_logic_vector(to_unsigned(240, 8)),
			7996 => std_logic_vector(to_unsigned(225, 8)),
			7997 => std_logic_vector(to_unsigned(166, 8)),
			7998 => std_logic_vector(to_unsigned(146, 8)),
			7999 => std_logic_vector(to_unsigned(64, 8)),
			8000 => std_logic_vector(to_unsigned(166, 8)),
			8001 => std_logic_vector(to_unsigned(52, 8)),
			8002 => std_logic_vector(to_unsigned(168, 8)),
			8003 => std_logic_vector(to_unsigned(206, 8)),
			8004 => std_logic_vector(to_unsigned(133, 8)),
			8005 => std_logic_vector(to_unsigned(48, 8)),
			8006 => std_logic_vector(to_unsigned(220, 8)),
			8007 => std_logic_vector(to_unsigned(6, 8)),
			8008 => std_logic_vector(to_unsigned(179, 8)),
			8009 => std_logic_vector(to_unsigned(137, 8)),
			8010 => std_logic_vector(to_unsigned(174, 8)),
			8011 => std_logic_vector(to_unsigned(67, 8)),
			8012 => std_logic_vector(to_unsigned(159, 8)),
			8013 => std_logic_vector(to_unsigned(187, 8)),
			8014 => std_logic_vector(to_unsigned(239, 8)),
			8015 => std_logic_vector(to_unsigned(236, 8)),
			8016 => std_logic_vector(to_unsigned(241, 8)),
			8017 => std_logic_vector(to_unsigned(225, 8)),
			8018 => std_logic_vector(to_unsigned(30, 8)),
			8019 => std_logic_vector(to_unsigned(142, 8)),
			8020 => std_logic_vector(to_unsigned(101, 8)),
			8021 => std_logic_vector(to_unsigned(233, 8)),
			8022 => std_logic_vector(to_unsigned(216, 8)),
			8023 => std_logic_vector(to_unsigned(132, 8)),
			8024 => std_logic_vector(to_unsigned(200, 8)),
			8025 => std_logic_vector(to_unsigned(63, 8)),
			8026 => std_logic_vector(to_unsigned(248, 8)),
			8027 => std_logic_vector(to_unsigned(152, 8)),
			8028 => std_logic_vector(to_unsigned(156, 8)),
			8029 => std_logic_vector(to_unsigned(119, 8)),
			8030 => std_logic_vector(to_unsigned(184, 8)),
			8031 => std_logic_vector(to_unsigned(232, 8)),
			8032 => std_logic_vector(to_unsigned(190, 8)),
			8033 => std_logic_vector(to_unsigned(165, 8)),
			8034 => std_logic_vector(to_unsigned(227, 8)),
			8035 => std_logic_vector(to_unsigned(0, 8)),
			8036 => std_logic_vector(to_unsigned(247, 8)),
			8037 => std_logic_vector(to_unsigned(15, 8)),
			8038 => std_logic_vector(to_unsigned(14, 8)),
			8039 => std_logic_vector(to_unsigned(174, 8)),
			8040 => std_logic_vector(to_unsigned(114, 8)),
			8041 => std_logic_vector(to_unsigned(252, 8)),
			8042 => std_logic_vector(to_unsigned(180, 8)),
			8043 => std_logic_vector(to_unsigned(39, 8)),
			8044 => std_logic_vector(to_unsigned(54, 8)),
			8045 => std_logic_vector(to_unsigned(9, 8)),
			8046 => std_logic_vector(to_unsigned(234, 8)),
			8047 => std_logic_vector(to_unsigned(0, 8)),
			8048 => std_logic_vector(to_unsigned(44, 8)),
			8049 => std_logic_vector(to_unsigned(247, 8)),
			8050 => std_logic_vector(to_unsigned(15, 8)),
			8051 => std_logic_vector(to_unsigned(83, 8)),
			8052 => std_logic_vector(to_unsigned(23, 8)),
			8053 => std_logic_vector(to_unsigned(203, 8)),
			8054 => std_logic_vector(to_unsigned(136, 8)),
			8055 => std_logic_vector(to_unsigned(153, 8)),
			8056 => std_logic_vector(to_unsigned(41, 8)),
			8057 => std_logic_vector(to_unsigned(39, 8)),
			8058 => std_logic_vector(to_unsigned(218, 8)),
			8059 => std_logic_vector(to_unsigned(74, 8)),
			8060 => std_logic_vector(to_unsigned(159, 8)),
			8061 => std_logic_vector(to_unsigned(65, 8)),
			8062 => std_logic_vector(to_unsigned(25, 8)),
			8063 => std_logic_vector(to_unsigned(169, 8)),
			8064 => std_logic_vector(to_unsigned(237, 8)),
			8065 => std_logic_vector(to_unsigned(106, 8)),
			8066 => std_logic_vector(to_unsigned(152, 8)),
			8067 => std_logic_vector(to_unsigned(21, 8)),
			8068 => std_logic_vector(to_unsigned(2, 8)),
			8069 => std_logic_vector(to_unsigned(154, 8)),
			8070 => std_logic_vector(to_unsigned(215, 8)),
			8071 => std_logic_vector(to_unsigned(125, 8)),
			8072 => std_logic_vector(to_unsigned(139, 8)),
			8073 => std_logic_vector(to_unsigned(95, 8)),
			8074 => std_logic_vector(to_unsigned(132, 8)),
			8075 => std_logic_vector(to_unsigned(88, 8)),
			8076 => std_logic_vector(to_unsigned(129, 8)),
			8077 => std_logic_vector(to_unsigned(36, 8)),
			8078 => std_logic_vector(to_unsigned(90, 8)),
			8079 => std_logic_vector(to_unsigned(125, 8)),
			8080 => std_logic_vector(to_unsigned(218, 8)),
			8081 => std_logic_vector(to_unsigned(41, 8)),
			8082 => std_logic_vector(to_unsigned(16, 8)),
			8083 => std_logic_vector(to_unsigned(214, 8)),
			8084 => std_logic_vector(to_unsigned(168, 8)),
			8085 => std_logic_vector(to_unsigned(122, 8)),
			8086 => std_logic_vector(to_unsigned(155, 8)),
			8087 => std_logic_vector(to_unsigned(94, 8)),
			8088 => std_logic_vector(to_unsigned(173, 8)),
			8089 => std_logic_vector(to_unsigned(6, 8)),
			8090 => std_logic_vector(to_unsigned(12, 8)),
			8091 => std_logic_vector(to_unsigned(8, 8)),
			8092 => std_logic_vector(to_unsigned(175, 8)),
			8093 => std_logic_vector(to_unsigned(34, 8)),
			8094 => std_logic_vector(to_unsigned(82, 8)),
			8095 => std_logic_vector(to_unsigned(89, 8)),
			8096 => std_logic_vector(to_unsigned(190, 8)),
			8097 => std_logic_vector(to_unsigned(135, 8)),
			8098 => std_logic_vector(to_unsigned(82, 8)),
			8099 => std_logic_vector(to_unsigned(253, 8)),
			8100 => std_logic_vector(to_unsigned(112, 8)),
			8101 => std_logic_vector(to_unsigned(104, 8)),
			8102 => std_logic_vector(to_unsigned(116, 8)),
			8103 => std_logic_vector(to_unsigned(111, 8)),
			8104 => std_logic_vector(to_unsigned(25, 8)),
			8105 => std_logic_vector(to_unsigned(68, 8)),
			8106 => std_logic_vector(to_unsigned(110, 8)),
			8107 => std_logic_vector(to_unsigned(219, 8)),
			8108 => std_logic_vector(to_unsigned(99, 8)),
			8109 => std_logic_vector(to_unsigned(105, 8)),
			8110 => std_logic_vector(to_unsigned(118, 8)),
			8111 => std_logic_vector(to_unsigned(223, 8)),
			8112 => std_logic_vector(to_unsigned(135, 8)),
			8113 => std_logic_vector(to_unsigned(45, 8)),
			8114 => std_logic_vector(to_unsigned(152, 8)),
			8115 => std_logic_vector(to_unsigned(200, 8)),
			8116 => std_logic_vector(to_unsigned(19, 8)),
			8117 => std_logic_vector(to_unsigned(209, 8)),
			8118 => std_logic_vector(to_unsigned(128, 8)),
			8119 => std_logic_vector(to_unsigned(162, 8)),
			8120 => std_logic_vector(to_unsigned(44, 8)),
			8121 => std_logic_vector(to_unsigned(52, 8)),
			8122 => std_logic_vector(to_unsigned(57, 8)),
			8123 => std_logic_vector(to_unsigned(75, 8)),
			8124 => std_logic_vector(to_unsigned(73, 8)),
			8125 => std_logic_vector(to_unsigned(235, 8)),
			8126 => std_logic_vector(to_unsigned(241, 8)),
			8127 => std_logic_vector(to_unsigned(245, 8)),
			8128 => std_logic_vector(to_unsigned(47, 8)),
			8129 => std_logic_vector(to_unsigned(50, 8)),
			8130 => std_logic_vector(to_unsigned(188, 8)),
			8131 => std_logic_vector(to_unsigned(187, 8)),
			8132 => std_logic_vector(to_unsigned(165, 8)),
			8133 => std_logic_vector(to_unsigned(36, 8)),
			8134 => std_logic_vector(to_unsigned(71, 8)),
			8135 => std_logic_vector(to_unsigned(193, 8)),
			8136 => std_logic_vector(to_unsigned(190, 8)),
			8137 => std_logic_vector(to_unsigned(108, 8)),
			8138 => std_logic_vector(to_unsigned(94, 8)),
			8139 => std_logic_vector(to_unsigned(24, 8)),
			8140 => std_logic_vector(to_unsigned(120, 8)),
			8141 => std_logic_vector(to_unsigned(29, 8)),
			8142 => std_logic_vector(to_unsigned(75, 8)),
			8143 => std_logic_vector(to_unsigned(10, 8)),
			8144 => std_logic_vector(to_unsigned(114, 8)),
			8145 => std_logic_vector(to_unsigned(167, 8)),
			8146 => std_logic_vector(to_unsigned(133, 8)),
			8147 => std_logic_vector(to_unsigned(45, 8)),
			8148 => std_logic_vector(to_unsigned(133, 8)),
			8149 => std_logic_vector(to_unsigned(50, 8)),
			8150 => std_logic_vector(to_unsigned(76, 8)),
			8151 => std_logic_vector(to_unsigned(54, 8)),
			8152 => std_logic_vector(to_unsigned(172, 8)),
			8153 => std_logic_vector(to_unsigned(174, 8)),
			8154 => std_logic_vector(to_unsigned(117, 8)),
			8155 => std_logic_vector(to_unsigned(165, 8)),
			8156 => std_logic_vector(to_unsigned(143, 8)),
			8157 => std_logic_vector(to_unsigned(184, 8)),
			8158 => std_logic_vector(to_unsigned(140, 8)),
			8159 => std_logic_vector(to_unsigned(191, 8)),
			8160 => std_logic_vector(to_unsigned(200, 8)),
			8161 => std_logic_vector(to_unsigned(177, 8)),
			8162 => std_logic_vector(to_unsigned(3, 8)),
			8163 => std_logic_vector(to_unsigned(51, 8)),
			8164 => std_logic_vector(to_unsigned(192, 8)),
			8165 => std_logic_vector(to_unsigned(86, 8)),
			8166 => std_logic_vector(to_unsigned(8, 8)),
			8167 => std_logic_vector(to_unsigned(11, 8)),
			8168 => std_logic_vector(to_unsigned(108, 8)),
			8169 => std_logic_vector(to_unsigned(183, 8)),
			8170 => std_logic_vector(to_unsigned(12, 8)),
			8171 => std_logic_vector(to_unsigned(11, 8)),
			8172 => std_logic_vector(to_unsigned(204, 8)),
			8173 => std_logic_vector(to_unsigned(68, 8)),
			8174 => std_logic_vector(to_unsigned(223, 8)),
			8175 => std_logic_vector(to_unsigned(95, 8)),
			8176 => std_logic_vector(to_unsigned(76, 8)),
			8177 => std_logic_vector(to_unsigned(172, 8)),
			8178 => std_logic_vector(to_unsigned(2, 8)),
			8179 => std_logic_vector(to_unsigned(157, 8)),
			8180 => std_logic_vector(to_unsigned(97, 8)),
			8181 => std_logic_vector(to_unsigned(77, 8)),
			8182 => std_logic_vector(to_unsigned(151, 8)),
			8183 => std_logic_vector(to_unsigned(173, 8)),
			8184 => std_logic_vector(to_unsigned(60, 8)),
			8185 => std_logic_vector(to_unsigned(171, 8)),
			8186 => std_logic_vector(to_unsigned(8, 8)),
			8187 => std_logic_vector(to_unsigned(125, 8)),
			8188 => std_logic_vector(to_unsigned(182, 8)),
			8189 => std_logic_vector(to_unsigned(5, 8)),
			8190 => std_logic_vector(to_unsigned(153, 8)),
			8191 => std_logic_vector(to_unsigned(37, 8)),
			8192 => std_logic_vector(to_unsigned(79, 8)),
			8193 => std_logic_vector(to_unsigned(120, 8)),
			8194 => std_logic_vector(to_unsigned(28, 8)),
			8195 => std_logic_vector(to_unsigned(156, 8)),
			8196 => std_logic_vector(to_unsigned(242, 8)),
			8197 => std_logic_vector(to_unsigned(6, 8)),
			8198 => std_logic_vector(to_unsigned(178, 8)),
			8199 => std_logic_vector(to_unsigned(7, 8)),
			8200 => std_logic_vector(to_unsigned(230, 8)),
			8201 => std_logic_vector(to_unsigned(82, 8)),
			8202 => std_logic_vector(to_unsigned(161, 8)),
			8203 => std_logic_vector(to_unsigned(186, 8)),
			8204 => std_logic_vector(to_unsigned(124, 8)),
			8205 => std_logic_vector(to_unsigned(210, 8)),
			8206 => std_logic_vector(to_unsigned(142, 8)),
			8207 => std_logic_vector(to_unsigned(203, 8)),
			8208 => std_logic_vector(to_unsigned(50, 8)),
			8209 => std_logic_vector(to_unsigned(142, 8)),
			8210 => std_logic_vector(to_unsigned(81, 8)),
			8211 => std_logic_vector(to_unsigned(145, 8)),
			8212 => std_logic_vector(to_unsigned(157, 8)),
			8213 => std_logic_vector(to_unsigned(192, 8)),
			8214 => std_logic_vector(to_unsigned(226, 8)),
			8215 => std_logic_vector(to_unsigned(88, 8)),
			8216 => std_logic_vector(to_unsigned(10, 8)),
			8217 => std_logic_vector(to_unsigned(110, 8)),
			8218 => std_logic_vector(to_unsigned(47, 8)),
			8219 => std_logic_vector(to_unsigned(62, 8)),
			8220 => std_logic_vector(to_unsigned(5, 8)),
			8221 => std_logic_vector(to_unsigned(136, 8)),
			8222 => std_logic_vector(to_unsigned(186, 8)),
			8223 => std_logic_vector(to_unsigned(109, 8)),
			8224 => std_logic_vector(to_unsigned(83, 8)),
			8225 => std_logic_vector(to_unsigned(120, 8)),
			8226 => std_logic_vector(to_unsigned(55, 8)),
			8227 => std_logic_vector(to_unsigned(100, 8)),
			8228 => std_logic_vector(to_unsigned(24, 8)),
			8229 => std_logic_vector(to_unsigned(234, 8)),
			8230 => std_logic_vector(to_unsigned(197, 8)),
			8231 => std_logic_vector(to_unsigned(9, 8)),
			8232 => std_logic_vector(to_unsigned(197, 8)),
			8233 => std_logic_vector(to_unsigned(162, 8)),
			8234 => std_logic_vector(to_unsigned(237, 8)),
			8235 => std_logic_vector(to_unsigned(108, 8)),
			8236 => std_logic_vector(to_unsigned(196, 8)),
			8237 => std_logic_vector(to_unsigned(134, 8)),
			8238 => std_logic_vector(to_unsigned(245, 8)),
			8239 => std_logic_vector(to_unsigned(25, 8)),
			8240 => std_logic_vector(to_unsigned(93, 8)),
			8241 => std_logic_vector(to_unsigned(1, 8)),
			8242 => std_logic_vector(to_unsigned(223, 8)),
			8243 => std_logic_vector(to_unsigned(125, 8)),
			8244 => std_logic_vector(to_unsigned(120, 8)),
			8245 => std_logic_vector(to_unsigned(228, 8)),
			8246 => std_logic_vector(to_unsigned(226, 8)),
			8247 => std_logic_vector(to_unsigned(122, 8)),
			8248 => std_logic_vector(to_unsigned(47, 8)),
			8249 => std_logic_vector(to_unsigned(101, 8)),
			8250 => std_logic_vector(to_unsigned(225, 8)),
			8251 => std_logic_vector(to_unsigned(228, 8)),
			8252 => std_logic_vector(to_unsigned(171, 8)),
			8253 => std_logic_vector(to_unsigned(83, 8)),
			8254 => std_logic_vector(to_unsigned(117, 8)),
			8255 => std_logic_vector(to_unsigned(208, 8)),
			8256 => std_logic_vector(to_unsigned(29, 8)),
			8257 => std_logic_vector(to_unsigned(192, 8)),
			8258 => std_logic_vector(to_unsigned(209, 8)),
			8259 => std_logic_vector(to_unsigned(217, 8)),
			8260 => std_logic_vector(to_unsigned(14, 8)),
			8261 => std_logic_vector(to_unsigned(207, 8)),
			8262 => std_logic_vector(to_unsigned(75, 8)),
			8263 => std_logic_vector(to_unsigned(71, 8)),
			8264 => std_logic_vector(to_unsigned(155, 8)),
			8265 => std_logic_vector(to_unsigned(230, 8)),
			8266 => std_logic_vector(to_unsigned(252, 8)),
			8267 => std_logic_vector(to_unsigned(14, 8)),
			8268 => std_logic_vector(to_unsigned(7, 8)),
			8269 => std_logic_vector(to_unsigned(118, 8)),
			8270 => std_logic_vector(to_unsigned(211, 8)),
			8271 => std_logic_vector(to_unsigned(37, 8)),
			8272 => std_logic_vector(to_unsigned(62, 8)),
			8273 => std_logic_vector(to_unsigned(214, 8)),
			8274 => std_logic_vector(to_unsigned(186, 8)),
			8275 => std_logic_vector(to_unsigned(242, 8)),
			8276 => std_logic_vector(to_unsigned(138, 8)),
			8277 => std_logic_vector(to_unsigned(3, 8)),
			8278 => std_logic_vector(to_unsigned(160, 8)),
			8279 => std_logic_vector(to_unsigned(97, 8)),
			8280 => std_logic_vector(to_unsigned(78, 8)),
			8281 => std_logic_vector(to_unsigned(198, 8)),
			8282 => std_logic_vector(to_unsigned(231, 8)),
			8283 => std_logic_vector(to_unsigned(4, 8)),
			8284 => std_logic_vector(to_unsigned(72, 8)),
			8285 => std_logic_vector(to_unsigned(199, 8)),
			8286 => std_logic_vector(to_unsigned(30, 8)),
			8287 => std_logic_vector(to_unsigned(132, 8)),
			8288 => std_logic_vector(to_unsigned(246, 8)),
			8289 => std_logic_vector(to_unsigned(115, 8)),
			8290 => std_logic_vector(to_unsigned(6, 8)),
			8291 => std_logic_vector(to_unsigned(213, 8)),
			8292 => std_logic_vector(to_unsigned(234, 8)),
			8293 => std_logic_vector(to_unsigned(153, 8)),
			8294 => std_logic_vector(to_unsigned(108, 8)),
			8295 => std_logic_vector(to_unsigned(207, 8)),
			8296 => std_logic_vector(to_unsigned(101, 8)),
			8297 => std_logic_vector(to_unsigned(181, 8)),
			8298 => std_logic_vector(to_unsigned(76, 8)),
			8299 => std_logic_vector(to_unsigned(94, 8)),
			8300 => std_logic_vector(to_unsigned(38, 8)),
			8301 => std_logic_vector(to_unsigned(66, 8)),
			8302 => std_logic_vector(to_unsigned(231, 8)),
			8303 => std_logic_vector(to_unsigned(102, 8)),
			8304 => std_logic_vector(to_unsigned(228, 8)),
			8305 => std_logic_vector(to_unsigned(177, 8)),
			8306 => std_logic_vector(to_unsigned(80, 8)),
			8307 => std_logic_vector(to_unsigned(170, 8)),
			8308 => std_logic_vector(to_unsigned(185, 8)),
			8309 => std_logic_vector(to_unsigned(22, 8)),
			8310 => std_logic_vector(to_unsigned(61, 8)),
			8311 => std_logic_vector(to_unsigned(242, 8)),
			8312 => std_logic_vector(to_unsigned(57, 8)),
			8313 => std_logic_vector(to_unsigned(203, 8)),
			8314 => std_logic_vector(to_unsigned(229, 8)),
			8315 => std_logic_vector(to_unsigned(68, 8)),
			8316 => std_logic_vector(to_unsigned(24, 8)),
			8317 => std_logic_vector(to_unsigned(62, 8)),
			8318 => std_logic_vector(to_unsigned(212, 8)),
			8319 => std_logic_vector(to_unsigned(190, 8)),
			8320 => std_logic_vector(to_unsigned(108, 8)),
			8321 => std_logic_vector(to_unsigned(38, 8)),
			8322 => std_logic_vector(to_unsigned(188, 8)),
			8323 => std_logic_vector(to_unsigned(97, 8)),
			8324 => std_logic_vector(to_unsigned(173, 8)),
			8325 => std_logic_vector(to_unsigned(64, 8)),
			8326 => std_logic_vector(to_unsigned(211, 8)),
			8327 => std_logic_vector(to_unsigned(194, 8)),
			8328 => std_logic_vector(to_unsigned(149, 8)),
			8329 => std_logic_vector(to_unsigned(7, 8)),
			8330 => std_logic_vector(to_unsigned(91, 8)),
			8331 => std_logic_vector(to_unsigned(229, 8)),
			8332 => std_logic_vector(to_unsigned(95, 8)),
			8333 => std_logic_vector(to_unsigned(48, 8)),
			8334 => std_logic_vector(to_unsigned(245, 8)),
			8335 => std_logic_vector(to_unsigned(246, 8)),
			8336 => std_logic_vector(to_unsigned(177, 8)),
			8337 => std_logic_vector(to_unsigned(39, 8)),
			8338 => std_logic_vector(to_unsigned(243, 8)),
			8339 => std_logic_vector(to_unsigned(249, 8)),
			8340 => std_logic_vector(to_unsigned(56, 8)),
			8341 => std_logic_vector(to_unsigned(230, 8)),
			8342 => std_logic_vector(to_unsigned(46, 8)),
			8343 => std_logic_vector(to_unsigned(94, 8)),
			8344 => std_logic_vector(to_unsigned(172, 8)),
			8345 => std_logic_vector(to_unsigned(48, 8)),
			8346 => std_logic_vector(to_unsigned(29, 8)),
			8347 => std_logic_vector(to_unsigned(217, 8)),
			8348 => std_logic_vector(to_unsigned(114, 8)),
			8349 => std_logic_vector(to_unsigned(75, 8)),
			8350 => std_logic_vector(to_unsigned(199, 8)),
			8351 => std_logic_vector(to_unsigned(231, 8)),
			8352 => std_logic_vector(to_unsigned(20, 8)),
			8353 => std_logic_vector(to_unsigned(223, 8)),
			8354 => std_logic_vector(to_unsigned(18, 8)),
			8355 => std_logic_vector(to_unsigned(197, 8)),
			8356 => std_logic_vector(to_unsigned(98, 8)),
			8357 => std_logic_vector(to_unsigned(113, 8)),
			8358 => std_logic_vector(to_unsigned(125, 8)),
			8359 => std_logic_vector(to_unsigned(9, 8)),
			8360 => std_logic_vector(to_unsigned(247, 8)),
			8361 => std_logic_vector(to_unsigned(96, 8)),
			8362 => std_logic_vector(to_unsigned(214, 8)),
			8363 => std_logic_vector(to_unsigned(15, 8)),
			8364 => std_logic_vector(to_unsigned(149, 8)),
			8365 => std_logic_vector(to_unsigned(238, 8)),
			8366 => std_logic_vector(to_unsigned(203, 8)),
			8367 => std_logic_vector(to_unsigned(237, 8)),
			8368 => std_logic_vector(to_unsigned(6, 8)),
			8369 => std_logic_vector(to_unsigned(240, 8)),
			8370 => std_logic_vector(to_unsigned(168, 8)),
			8371 => std_logic_vector(to_unsigned(201, 8)),
			8372 => std_logic_vector(to_unsigned(232, 8)),
			8373 => std_logic_vector(to_unsigned(159, 8)),
			8374 => std_logic_vector(to_unsigned(190, 8)),
			8375 => std_logic_vector(to_unsigned(51, 8)),
			8376 => std_logic_vector(to_unsigned(54, 8)),
			8377 => std_logic_vector(to_unsigned(150, 8)),
			8378 => std_logic_vector(to_unsigned(59, 8)),
			8379 => std_logic_vector(to_unsigned(8, 8)),
			8380 => std_logic_vector(to_unsigned(23, 8)),
			8381 => std_logic_vector(to_unsigned(42, 8)),
			8382 => std_logic_vector(to_unsigned(124, 8)),
			8383 => std_logic_vector(to_unsigned(157, 8)),
			8384 => std_logic_vector(to_unsigned(155, 8)),
			8385 => std_logic_vector(to_unsigned(189, 8)),
			8386 => std_logic_vector(to_unsigned(245, 8)),
			8387 => std_logic_vector(to_unsigned(32, 8)),
			8388 => std_logic_vector(to_unsigned(131, 8)),
			8389 => std_logic_vector(to_unsigned(155, 8)),
			8390 => std_logic_vector(to_unsigned(61, 8)),
			8391 => std_logic_vector(to_unsigned(97, 8)),
			8392 => std_logic_vector(to_unsigned(173, 8)),
			8393 => std_logic_vector(to_unsigned(55, 8)),
			8394 => std_logic_vector(to_unsigned(69, 8)),
			8395 => std_logic_vector(to_unsigned(57, 8)),
			8396 => std_logic_vector(to_unsigned(174, 8)),
			8397 => std_logic_vector(to_unsigned(6, 8)),
			8398 => std_logic_vector(to_unsigned(212, 8)),
			8399 => std_logic_vector(to_unsigned(234, 8)),
			8400 => std_logic_vector(to_unsigned(241, 8)),
			8401 => std_logic_vector(to_unsigned(3, 8)),
			8402 => std_logic_vector(to_unsigned(185, 8)),
			8403 => std_logic_vector(to_unsigned(168, 8)),
			8404 => std_logic_vector(to_unsigned(57, 8)),
			8405 => std_logic_vector(to_unsigned(131, 8)),
			8406 => std_logic_vector(to_unsigned(13, 8)),
			8407 => std_logic_vector(to_unsigned(164, 8)),
			8408 => std_logic_vector(to_unsigned(13, 8)),
			8409 => std_logic_vector(to_unsigned(101, 8)),
			8410 => std_logic_vector(to_unsigned(219, 8)),
			8411 => std_logic_vector(to_unsigned(81, 8)),
			8412 => std_logic_vector(to_unsigned(231, 8)),
			8413 => std_logic_vector(to_unsigned(122, 8)),
			8414 => std_logic_vector(to_unsigned(73, 8)),
			8415 => std_logic_vector(to_unsigned(132, 8)),
			8416 => std_logic_vector(to_unsigned(141, 8)),
			8417 => std_logic_vector(to_unsigned(207, 8)),
			8418 => std_logic_vector(to_unsigned(143, 8)),
			8419 => std_logic_vector(to_unsigned(151, 8)),
			8420 => std_logic_vector(to_unsigned(70, 8)),
			8421 => std_logic_vector(to_unsigned(247, 8)),
			8422 => std_logic_vector(to_unsigned(9, 8)),
			8423 => std_logic_vector(to_unsigned(229, 8)),
			8424 => std_logic_vector(to_unsigned(90, 8)),
			8425 => std_logic_vector(to_unsigned(134, 8)),
			8426 => std_logic_vector(to_unsigned(196, 8)),
			8427 => std_logic_vector(to_unsigned(6, 8)),
			8428 => std_logic_vector(to_unsigned(146, 8)),
			8429 => std_logic_vector(to_unsigned(140, 8)),
			8430 => std_logic_vector(to_unsigned(58, 8)),
			8431 => std_logic_vector(to_unsigned(78, 8)),
			8432 => std_logic_vector(to_unsigned(42, 8)),
			8433 => std_logic_vector(to_unsigned(53, 8)),
			8434 => std_logic_vector(to_unsigned(43, 8)),
			8435 => std_logic_vector(to_unsigned(38, 8)),
			8436 => std_logic_vector(to_unsigned(87, 8)),
			8437 => std_logic_vector(to_unsigned(246, 8)),
			8438 => std_logic_vector(to_unsigned(88, 8)),
			8439 => std_logic_vector(to_unsigned(169, 8)),
			8440 => std_logic_vector(to_unsigned(158, 8)),
			8441 => std_logic_vector(to_unsigned(103, 8)),
			8442 => std_logic_vector(to_unsigned(50, 8)),
			8443 => std_logic_vector(to_unsigned(31, 8)),
			8444 => std_logic_vector(to_unsigned(120, 8)),
			8445 => std_logic_vector(to_unsigned(46, 8)),
			8446 => std_logic_vector(to_unsigned(67, 8)),
			8447 => std_logic_vector(to_unsigned(48, 8)),
			8448 => std_logic_vector(to_unsigned(1, 8)),
			8449 => std_logic_vector(to_unsigned(164, 8)),
			8450 => std_logic_vector(to_unsigned(76, 8)),
			8451 => std_logic_vector(to_unsigned(179, 8)),
			8452 => std_logic_vector(to_unsigned(106, 8)),
			8453 => std_logic_vector(to_unsigned(107, 8)),
			8454 => std_logic_vector(to_unsigned(153, 8)),
			8455 => std_logic_vector(to_unsigned(10, 8)),
			8456 => std_logic_vector(to_unsigned(29, 8)),
			8457 => std_logic_vector(to_unsigned(200, 8)),
			8458 => std_logic_vector(to_unsigned(221, 8)),
			8459 => std_logic_vector(to_unsigned(219, 8)),
			8460 => std_logic_vector(to_unsigned(32, 8)),
			8461 => std_logic_vector(to_unsigned(7, 8)),
			8462 => std_logic_vector(to_unsigned(107, 8)),
			8463 => std_logic_vector(to_unsigned(20, 8)),
			8464 => std_logic_vector(to_unsigned(117, 8)),
			8465 => std_logic_vector(to_unsigned(74, 8)),
			8466 => std_logic_vector(to_unsigned(154, 8)),
			8467 => std_logic_vector(to_unsigned(66, 8)),
			8468 => std_logic_vector(to_unsigned(126, 8)),
			8469 => std_logic_vector(to_unsigned(131, 8)),
			8470 => std_logic_vector(to_unsigned(33, 8)),
			8471 => std_logic_vector(to_unsigned(127, 8)),
			8472 => std_logic_vector(to_unsigned(233, 8)),
			8473 => std_logic_vector(to_unsigned(104, 8)),
			8474 => std_logic_vector(to_unsigned(153, 8)),
			8475 => std_logic_vector(to_unsigned(110, 8)),
			8476 => std_logic_vector(to_unsigned(253, 8)),
			8477 => std_logic_vector(to_unsigned(43, 8)),
			8478 => std_logic_vector(to_unsigned(172, 8)),
			8479 => std_logic_vector(to_unsigned(175, 8)),
			8480 => std_logic_vector(to_unsigned(117, 8)),
			8481 => std_logic_vector(to_unsigned(163, 8)),
			8482 => std_logic_vector(to_unsigned(8, 8)),
			8483 => std_logic_vector(to_unsigned(104, 8)),
			8484 => std_logic_vector(to_unsigned(118, 8)),
			8485 => std_logic_vector(to_unsigned(41, 8)),
			8486 => std_logic_vector(to_unsigned(202, 8)),
			8487 => std_logic_vector(to_unsigned(123, 8)),
			8488 => std_logic_vector(to_unsigned(98, 8)),
			8489 => std_logic_vector(to_unsigned(13, 8)),
			8490 => std_logic_vector(to_unsigned(123, 8)),
			8491 => std_logic_vector(to_unsigned(28, 8)),
			8492 => std_logic_vector(to_unsigned(129, 8)),
			8493 => std_logic_vector(to_unsigned(204, 8)),
			8494 => std_logic_vector(to_unsigned(23, 8)),
			8495 => std_logic_vector(to_unsigned(71, 8)),
			8496 => std_logic_vector(to_unsigned(198, 8)),
			8497 => std_logic_vector(to_unsigned(12, 8)),
			8498 => std_logic_vector(to_unsigned(147, 8)),
			8499 => std_logic_vector(to_unsigned(238, 8)),
			8500 => std_logic_vector(to_unsigned(114, 8)),
			8501 => std_logic_vector(to_unsigned(20, 8)),
			8502 => std_logic_vector(to_unsigned(213, 8)),
			8503 => std_logic_vector(to_unsigned(254, 8)),
			8504 => std_logic_vector(to_unsigned(199, 8)),
			8505 => std_logic_vector(to_unsigned(155, 8)),
			8506 => std_logic_vector(to_unsigned(34, 8)),
			8507 => std_logic_vector(to_unsigned(128, 8)),
			8508 => std_logic_vector(to_unsigned(99, 8)),
			8509 => std_logic_vector(to_unsigned(4, 8)),
			8510 => std_logic_vector(to_unsigned(155, 8)),
			8511 => std_logic_vector(to_unsigned(36, 8)),
			8512 => std_logic_vector(to_unsigned(43, 8)),
			8513 => std_logic_vector(to_unsigned(210, 8)),
			8514 => std_logic_vector(to_unsigned(93, 8)),
			8515 => std_logic_vector(to_unsigned(174, 8)),
			8516 => std_logic_vector(to_unsigned(248, 8)),
			8517 => std_logic_vector(to_unsigned(26, 8)),
			8518 => std_logic_vector(to_unsigned(68, 8)),
			8519 => std_logic_vector(to_unsigned(183, 8)),
			8520 => std_logic_vector(to_unsigned(209, 8)),
			8521 => std_logic_vector(to_unsigned(82, 8)),
			8522 => std_logic_vector(to_unsigned(80, 8)),
			8523 => std_logic_vector(to_unsigned(200, 8)),
			8524 => std_logic_vector(to_unsigned(63, 8)),
			8525 => std_logic_vector(to_unsigned(107, 8)),
			8526 => std_logic_vector(to_unsigned(36, 8)),
			8527 => std_logic_vector(to_unsigned(67, 8)),
			8528 => std_logic_vector(to_unsigned(70, 8)),
			8529 => std_logic_vector(to_unsigned(122, 8)),
			8530 => std_logic_vector(to_unsigned(57, 8)),
			8531 => std_logic_vector(to_unsigned(206, 8)),
			8532 => std_logic_vector(to_unsigned(1, 8)),
			8533 => std_logic_vector(to_unsigned(143, 8)),
			8534 => std_logic_vector(to_unsigned(228, 8)),
			8535 => std_logic_vector(to_unsigned(137, 8)),
			8536 => std_logic_vector(to_unsigned(56, 8)),
			8537 => std_logic_vector(to_unsigned(163, 8)),
			8538 => std_logic_vector(to_unsigned(119, 8)),
			8539 => std_logic_vector(to_unsigned(129, 8)),
			8540 => std_logic_vector(to_unsigned(196, 8)),
			8541 => std_logic_vector(to_unsigned(76, 8)),
			8542 => std_logic_vector(to_unsigned(53, 8)),
			8543 => std_logic_vector(to_unsigned(245, 8)),
			8544 => std_logic_vector(to_unsigned(19, 8)),
			8545 => std_logic_vector(to_unsigned(178, 8)),
			8546 => std_logic_vector(to_unsigned(198, 8)),
			8547 => std_logic_vector(to_unsigned(246, 8)),
			8548 => std_logic_vector(to_unsigned(13, 8)),
			8549 => std_logic_vector(to_unsigned(20, 8)),
			8550 => std_logic_vector(to_unsigned(198, 8)),
			8551 => std_logic_vector(to_unsigned(147, 8)),
			8552 => std_logic_vector(to_unsigned(187, 8)),
			8553 => std_logic_vector(to_unsigned(239, 8)),
			8554 => std_logic_vector(to_unsigned(124, 8)),
			8555 => std_logic_vector(to_unsigned(131, 8)),
			8556 => std_logic_vector(to_unsigned(66, 8)),
			8557 => std_logic_vector(to_unsigned(130, 8)),
			8558 => std_logic_vector(to_unsigned(202, 8)),
			8559 => std_logic_vector(to_unsigned(98, 8)),
			8560 => std_logic_vector(to_unsigned(108, 8)),
			8561 => std_logic_vector(to_unsigned(83, 8)),
			8562 => std_logic_vector(to_unsigned(185, 8)),
			8563 => std_logic_vector(to_unsigned(148, 8)),
			8564 => std_logic_vector(to_unsigned(169, 8)),
			8565 => std_logic_vector(to_unsigned(35, 8)),
			8566 => std_logic_vector(to_unsigned(127, 8)),
			8567 => std_logic_vector(to_unsigned(71, 8)),
			8568 => std_logic_vector(to_unsigned(201, 8)),
			8569 => std_logic_vector(to_unsigned(12, 8)),
			8570 => std_logic_vector(to_unsigned(18, 8)),
			8571 => std_logic_vector(to_unsigned(12, 8)),
			8572 => std_logic_vector(to_unsigned(158, 8)),
			8573 => std_logic_vector(to_unsigned(175, 8)),
			8574 => std_logic_vector(to_unsigned(107, 8)),
			8575 => std_logic_vector(to_unsigned(187, 8)),
			8576 => std_logic_vector(to_unsigned(183, 8)),
			8577 => std_logic_vector(to_unsigned(204, 8)),
			8578 => std_logic_vector(to_unsigned(162, 8)),
			8579 => std_logic_vector(to_unsigned(220, 8)),
			8580 => std_logic_vector(to_unsigned(99, 8)),
			8581 => std_logic_vector(to_unsigned(221, 8)),
			8582 => std_logic_vector(to_unsigned(230, 8)),
			8583 => std_logic_vector(to_unsigned(135, 8)),
			8584 => std_logic_vector(to_unsigned(128, 8)),
			8585 => std_logic_vector(to_unsigned(1, 8)),
			8586 => std_logic_vector(to_unsigned(137, 8)),
			8587 => std_logic_vector(to_unsigned(70, 8)),
			8588 => std_logic_vector(to_unsigned(69, 8)),
			8589 => std_logic_vector(to_unsigned(51, 8)),
			8590 => std_logic_vector(to_unsigned(91, 8)),
			8591 => std_logic_vector(to_unsigned(156, 8)),
			8592 => std_logic_vector(to_unsigned(91, 8)),
			8593 => std_logic_vector(to_unsigned(112, 8)),
			8594 => std_logic_vector(to_unsigned(31, 8)),
			8595 => std_logic_vector(to_unsigned(25, 8)),
			8596 => std_logic_vector(to_unsigned(109, 8)),
			8597 => std_logic_vector(to_unsigned(183, 8)),
			8598 => std_logic_vector(to_unsigned(247, 8)),
			8599 => std_logic_vector(to_unsigned(7, 8)),
			8600 => std_logic_vector(to_unsigned(40, 8)),
			8601 => std_logic_vector(to_unsigned(206, 8)),
			8602 => std_logic_vector(to_unsigned(252, 8)),
			8603 => std_logic_vector(to_unsigned(205, 8)),
			8604 => std_logic_vector(to_unsigned(186, 8)),
			8605 => std_logic_vector(to_unsigned(148, 8)),
			8606 => std_logic_vector(to_unsigned(153, 8)),
			8607 => std_logic_vector(to_unsigned(130, 8)),
			8608 => std_logic_vector(to_unsigned(120, 8)),
			8609 => std_logic_vector(to_unsigned(115, 8)),
			8610 => std_logic_vector(to_unsigned(172, 8)),
			8611 => std_logic_vector(to_unsigned(137, 8)),
			8612 => std_logic_vector(to_unsigned(0, 8)),
			8613 => std_logic_vector(to_unsigned(175, 8)),
			8614 => std_logic_vector(to_unsigned(216, 8)),
			8615 => std_logic_vector(to_unsigned(150, 8)),
			8616 => std_logic_vector(to_unsigned(158, 8)),
			8617 => std_logic_vector(to_unsigned(75, 8)),
			8618 => std_logic_vector(to_unsigned(95, 8)),
			8619 => std_logic_vector(to_unsigned(8, 8)),
			8620 => std_logic_vector(to_unsigned(82, 8)),
			8621 => std_logic_vector(to_unsigned(15, 8)),
			8622 => std_logic_vector(to_unsigned(212, 8)),
			8623 => std_logic_vector(to_unsigned(38, 8)),
			8624 => std_logic_vector(to_unsigned(1, 8)),
			8625 => std_logic_vector(to_unsigned(12, 8)),
			8626 => std_logic_vector(to_unsigned(232, 8)),
			8627 => std_logic_vector(to_unsigned(139, 8)),
			8628 => std_logic_vector(to_unsigned(216, 8)),
			8629 => std_logic_vector(to_unsigned(220, 8)),
			8630 => std_logic_vector(to_unsigned(203, 8)),
			8631 => std_logic_vector(to_unsigned(17, 8)),
			8632 => std_logic_vector(to_unsigned(70, 8)),
			8633 => std_logic_vector(to_unsigned(193, 8)),
			8634 => std_logic_vector(to_unsigned(32, 8)),
			8635 => std_logic_vector(to_unsigned(187, 8)),
			8636 => std_logic_vector(to_unsigned(193, 8)),
			8637 => std_logic_vector(to_unsigned(75, 8)),
			8638 => std_logic_vector(to_unsigned(14, 8)),
			8639 => std_logic_vector(to_unsigned(107, 8)),
			8640 => std_logic_vector(to_unsigned(240, 8)),
			8641 => std_logic_vector(to_unsigned(188, 8)),
			8642 => std_logic_vector(to_unsigned(63, 8)),
			8643 => std_logic_vector(to_unsigned(205, 8)),
			8644 => std_logic_vector(to_unsigned(35, 8)),
			8645 => std_logic_vector(to_unsigned(236, 8)),
			8646 => std_logic_vector(to_unsigned(151, 8)),
			8647 => std_logic_vector(to_unsigned(55, 8)),
			8648 => std_logic_vector(to_unsigned(26, 8)),
			8649 => std_logic_vector(to_unsigned(57, 8)),
			8650 => std_logic_vector(to_unsigned(66, 8)),
			8651 => std_logic_vector(to_unsigned(216, 8)),
			8652 => std_logic_vector(to_unsigned(172, 8)),
			8653 => std_logic_vector(to_unsigned(196, 8)),
			8654 => std_logic_vector(to_unsigned(61, 8)),
			8655 => std_logic_vector(to_unsigned(102, 8)),
			8656 => std_logic_vector(to_unsigned(208, 8)),
			8657 => std_logic_vector(to_unsigned(181, 8)),
			8658 => std_logic_vector(to_unsigned(182, 8)),
			8659 => std_logic_vector(to_unsigned(183, 8)),
			8660 => std_logic_vector(to_unsigned(239, 8)),
			8661 => std_logic_vector(to_unsigned(13, 8)),
			8662 => std_logic_vector(to_unsigned(169, 8)),
			8663 => std_logic_vector(to_unsigned(49, 8)),
			8664 => std_logic_vector(to_unsigned(183, 8)),
			8665 => std_logic_vector(to_unsigned(203, 8)),
			8666 => std_logic_vector(to_unsigned(95, 8)),
			8667 => std_logic_vector(to_unsigned(139, 8)),
			8668 => std_logic_vector(to_unsigned(213, 8)),
			8669 => std_logic_vector(to_unsigned(156, 8)),
			8670 => std_logic_vector(to_unsigned(87, 8)),
			8671 => std_logic_vector(to_unsigned(154, 8)),
			8672 => std_logic_vector(to_unsigned(68, 8)),
			8673 => std_logic_vector(to_unsigned(137, 8)),
			8674 => std_logic_vector(to_unsigned(181, 8)),
			8675 => std_logic_vector(to_unsigned(212, 8)),
			8676 => std_logic_vector(to_unsigned(208, 8)),
			8677 => std_logic_vector(to_unsigned(209, 8)),
			8678 => std_logic_vector(to_unsigned(134, 8)),
			8679 => std_logic_vector(to_unsigned(186, 8)),
			8680 => std_logic_vector(to_unsigned(195, 8)),
			8681 => std_logic_vector(to_unsigned(236, 8)),
			8682 => std_logic_vector(to_unsigned(99, 8)),
			8683 => std_logic_vector(to_unsigned(131, 8)),
			8684 => std_logic_vector(to_unsigned(175, 8)),
			8685 => std_logic_vector(to_unsigned(112, 8)),
			8686 => std_logic_vector(to_unsigned(117, 8)),
			8687 => std_logic_vector(to_unsigned(120, 8)),
			8688 => std_logic_vector(to_unsigned(127, 8)),
			8689 => std_logic_vector(to_unsigned(177, 8)),
			8690 => std_logic_vector(to_unsigned(191, 8)),
			8691 => std_logic_vector(to_unsigned(63, 8)),
			8692 => std_logic_vector(to_unsigned(176, 8)),
			8693 => std_logic_vector(to_unsigned(246, 8)),
			8694 => std_logic_vector(to_unsigned(145, 8)),
			8695 => std_logic_vector(to_unsigned(31, 8)),
			8696 => std_logic_vector(to_unsigned(80, 8)),
			8697 => std_logic_vector(to_unsigned(148, 8)),
			8698 => std_logic_vector(to_unsigned(44, 8)),
			8699 => std_logic_vector(to_unsigned(142, 8)),
			8700 => std_logic_vector(to_unsigned(71, 8)),
			8701 => std_logic_vector(to_unsigned(40, 8)),
			8702 => std_logic_vector(to_unsigned(237, 8)),
			8703 => std_logic_vector(to_unsigned(4, 8)),
			8704 => std_logic_vector(to_unsigned(248, 8)),
			8705 => std_logic_vector(to_unsigned(227, 8)),
			8706 => std_logic_vector(to_unsigned(82, 8)),
			8707 => std_logic_vector(to_unsigned(218, 8)),
			8708 => std_logic_vector(to_unsigned(28, 8)),
			8709 => std_logic_vector(to_unsigned(143, 8)),
			8710 => std_logic_vector(to_unsigned(197, 8)),
			8711 => std_logic_vector(to_unsigned(42, 8)),
			8712 => std_logic_vector(to_unsigned(49, 8)),
			8713 => std_logic_vector(to_unsigned(29, 8)),
			8714 => std_logic_vector(to_unsigned(112, 8)),
			8715 => std_logic_vector(to_unsigned(36, 8)),
			8716 => std_logic_vector(to_unsigned(107, 8)),
			8717 => std_logic_vector(to_unsigned(250, 8)),
			8718 => std_logic_vector(to_unsigned(82, 8)),
			8719 => std_logic_vector(to_unsigned(62, 8)),
			8720 => std_logic_vector(to_unsigned(109, 8)),
			8721 => std_logic_vector(to_unsigned(208, 8)),
			8722 => std_logic_vector(to_unsigned(205, 8)),
			8723 => std_logic_vector(to_unsigned(161, 8)),
			8724 => std_logic_vector(to_unsigned(113, 8)),
			8725 => std_logic_vector(to_unsigned(180, 8)),
			8726 => std_logic_vector(to_unsigned(189, 8)),
			8727 => std_logic_vector(to_unsigned(232, 8)),
			8728 => std_logic_vector(to_unsigned(248, 8)),
			8729 => std_logic_vector(to_unsigned(175, 8)),
			8730 => std_logic_vector(to_unsigned(166, 8)),
			8731 => std_logic_vector(to_unsigned(102, 8)),
			8732 => std_logic_vector(to_unsigned(248, 8)),
			8733 => std_logic_vector(to_unsigned(69, 8)),
			8734 => std_logic_vector(to_unsigned(15, 8)),
			8735 => std_logic_vector(to_unsigned(144, 8)),
			8736 => std_logic_vector(to_unsigned(40, 8)),
			8737 => std_logic_vector(to_unsigned(68, 8)),
			8738 => std_logic_vector(to_unsigned(227, 8)),
			8739 => std_logic_vector(to_unsigned(254, 8)),
			8740 => std_logic_vector(to_unsigned(41, 8)),
			8741 => std_logic_vector(to_unsigned(126, 8)),
			8742 => std_logic_vector(to_unsigned(35, 8)),
			8743 => std_logic_vector(to_unsigned(146, 8)),
			8744 => std_logic_vector(to_unsigned(221, 8)),
			8745 => std_logic_vector(to_unsigned(35, 8)),
			8746 => std_logic_vector(to_unsigned(6, 8)),
			8747 => std_logic_vector(to_unsigned(196, 8)),
			8748 => std_logic_vector(to_unsigned(78, 8)),
			8749 => std_logic_vector(to_unsigned(72, 8)),
			8750 => std_logic_vector(to_unsigned(189, 8)),
			8751 => std_logic_vector(to_unsigned(220, 8)),
			8752 => std_logic_vector(to_unsigned(225, 8)),
			8753 => std_logic_vector(to_unsigned(192, 8)),
			8754 => std_logic_vector(to_unsigned(249, 8)),
			8755 => std_logic_vector(to_unsigned(156, 8)),
			8756 => std_logic_vector(to_unsigned(198, 8)),
			8757 => std_logic_vector(to_unsigned(152, 8)),
			8758 => std_logic_vector(to_unsigned(106, 8)),
			8759 => std_logic_vector(to_unsigned(53, 8)),
			8760 => std_logic_vector(to_unsigned(169, 8)),
			8761 => std_logic_vector(to_unsigned(221, 8)),
			8762 => std_logic_vector(to_unsigned(244, 8)),
			8763 => std_logic_vector(to_unsigned(154, 8)),
			8764 => std_logic_vector(to_unsigned(163, 8)),
			8765 => std_logic_vector(to_unsigned(71, 8)),
			8766 => std_logic_vector(to_unsigned(196, 8)),
			8767 => std_logic_vector(to_unsigned(8, 8)),
			8768 => std_logic_vector(to_unsigned(73, 8)),
			8769 => std_logic_vector(to_unsigned(176, 8)),
			8770 => std_logic_vector(to_unsigned(227, 8)),
			8771 => std_logic_vector(to_unsigned(176, 8)),
			8772 => std_logic_vector(to_unsigned(165, 8)),
			8773 => std_logic_vector(to_unsigned(47, 8)),
			8774 => std_logic_vector(to_unsigned(218, 8)),
			8775 => std_logic_vector(to_unsigned(25, 8)),
			8776 => std_logic_vector(to_unsigned(184, 8)),
			8777 => std_logic_vector(to_unsigned(255, 8)),
			8778 => std_logic_vector(to_unsigned(72, 8)),
			8779 => std_logic_vector(to_unsigned(154, 8)),
			8780 => std_logic_vector(to_unsigned(59, 8)),
			8781 => std_logic_vector(to_unsigned(185, 8)),
			8782 => std_logic_vector(to_unsigned(20, 8)),
			8783 => std_logic_vector(to_unsigned(38, 8)),
			8784 => std_logic_vector(to_unsigned(50, 8)),
			8785 => std_logic_vector(to_unsigned(61, 8)),
			8786 => std_logic_vector(to_unsigned(114, 8)),
			8787 => std_logic_vector(to_unsigned(12, 8)),
			8788 => std_logic_vector(to_unsigned(114, 8)),
			8789 => std_logic_vector(to_unsigned(110, 8)),
			8790 => std_logic_vector(to_unsigned(93, 8)),
			8791 => std_logic_vector(to_unsigned(101, 8)),
			8792 => std_logic_vector(to_unsigned(130, 8)),
			8793 => std_logic_vector(to_unsigned(167, 8)),
			8794 => std_logic_vector(to_unsigned(151, 8)),
			8795 => std_logic_vector(to_unsigned(201, 8)),
			8796 => std_logic_vector(to_unsigned(24, 8)),
			8797 => std_logic_vector(to_unsigned(166, 8)),
			8798 => std_logic_vector(to_unsigned(23, 8)),
			8799 => std_logic_vector(to_unsigned(93, 8)),
			8800 => std_logic_vector(to_unsigned(203, 8)),
			8801 => std_logic_vector(to_unsigned(115, 8)),
			8802 => std_logic_vector(to_unsigned(139, 8)),
			8803 => std_logic_vector(to_unsigned(88, 8)),
			8804 => std_logic_vector(to_unsigned(136, 8)),
			8805 => std_logic_vector(to_unsigned(9, 8)),
			8806 => std_logic_vector(to_unsigned(20, 8)),
			8807 => std_logic_vector(to_unsigned(1, 8)),
			8808 => std_logic_vector(to_unsigned(58, 8)),
			8809 => std_logic_vector(to_unsigned(14, 8)),
			8810 => std_logic_vector(to_unsigned(106, 8)),
			8811 => std_logic_vector(to_unsigned(126, 8)),
			8812 => std_logic_vector(to_unsigned(97, 8)),
			8813 => std_logic_vector(to_unsigned(160, 8)),
			8814 => std_logic_vector(to_unsigned(97, 8)),
			8815 => std_logic_vector(to_unsigned(139, 8)),
			8816 => std_logic_vector(to_unsigned(220, 8)),
			8817 => std_logic_vector(to_unsigned(4, 8)),
			8818 => std_logic_vector(to_unsigned(123, 8)),
			8819 => std_logic_vector(to_unsigned(43, 8)),
			8820 => std_logic_vector(to_unsigned(145, 8)),
			8821 => std_logic_vector(to_unsigned(24, 8)),
			8822 => std_logic_vector(to_unsigned(95, 8)),
			8823 => std_logic_vector(to_unsigned(65, 8)),
			8824 => std_logic_vector(to_unsigned(1, 8)),
			8825 => std_logic_vector(to_unsigned(13, 8)),
			8826 => std_logic_vector(to_unsigned(74, 8)),
			8827 => std_logic_vector(to_unsigned(124, 8)),
			8828 => std_logic_vector(to_unsigned(12, 8)),
			8829 => std_logic_vector(to_unsigned(63, 8)),
			8830 => std_logic_vector(to_unsigned(112, 8)),
			8831 => std_logic_vector(to_unsigned(10, 8)),
			8832 => std_logic_vector(to_unsigned(233, 8)),
			8833 => std_logic_vector(to_unsigned(132, 8)),
			8834 => std_logic_vector(to_unsigned(240, 8)),
			8835 => std_logic_vector(to_unsigned(162, 8)),
			8836 => std_logic_vector(to_unsigned(64, 8)),
			8837 => std_logic_vector(to_unsigned(111, 8)),
			8838 => std_logic_vector(to_unsigned(154, 8)),
			8839 => std_logic_vector(to_unsigned(37, 8)),
			8840 => std_logic_vector(to_unsigned(233, 8)),
			8841 => std_logic_vector(to_unsigned(201, 8)),
			8842 => std_logic_vector(to_unsigned(124, 8)),
			8843 => std_logic_vector(to_unsigned(158, 8)),
			8844 => std_logic_vector(to_unsigned(55, 8)),
			8845 => std_logic_vector(to_unsigned(80, 8)),
			8846 => std_logic_vector(to_unsigned(246, 8)),
			8847 => std_logic_vector(to_unsigned(206, 8)),
			8848 => std_logic_vector(to_unsigned(55, 8)),
			8849 => std_logic_vector(to_unsigned(137, 8)),
			8850 => std_logic_vector(to_unsigned(109, 8)),
			8851 => std_logic_vector(to_unsigned(234, 8)),
			8852 => std_logic_vector(to_unsigned(131, 8)),
			8853 => std_logic_vector(to_unsigned(155, 8)),
			8854 => std_logic_vector(to_unsigned(56, 8)),
			8855 => std_logic_vector(to_unsigned(237, 8)),
			8856 => std_logic_vector(to_unsigned(216, 8)),
			8857 => std_logic_vector(to_unsigned(14, 8)),
			8858 => std_logic_vector(to_unsigned(155, 8)),
			8859 => std_logic_vector(to_unsigned(166, 8)),
			8860 => std_logic_vector(to_unsigned(172, 8)),
			8861 => std_logic_vector(to_unsigned(148, 8)),
			8862 => std_logic_vector(to_unsigned(50, 8)),
			8863 => std_logic_vector(to_unsigned(69, 8)),
			8864 => std_logic_vector(to_unsigned(186, 8)),
			8865 => std_logic_vector(to_unsigned(111, 8)),
			8866 => std_logic_vector(to_unsigned(188, 8)),
			8867 => std_logic_vector(to_unsigned(158, 8)),
			8868 => std_logic_vector(to_unsigned(149, 8)),
			8869 => std_logic_vector(to_unsigned(132, 8)),
			8870 => std_logic_vector(to_unsigned(137, 8)),
			8871 => std_logic_vector(to_unsigned(29, 8)),
			8872 => std_logic_vector(to_unsigned(31, 8)),
			8873 => std_logic_vector(to_unsigned(30, 8)),
			8874 => std_logic_vector(to_unsigned(53, 8)),
			8875 => std_logic_vector(to_unsigned(248, 8)),
			8876 => std_logic_vector(to_unsigned(137, 8)),
			8877 => std_logic_vector(to_unsigned(90, 8)),
			8878 => std_logic_vector(to_unsigned(58, 8)),
			8879 => std_logic_vector(to_unsigned(157, 8)),
			8880 => std_logic_vector(to_unsigned(156, 8)),
			8881 => std_logic_vector(to_unsigned(140, 8)),
			8882 => std_logic_vector(to_unsigned(112, 8)),
			8883 => std_logic_vector(to_unsigned(203, 8)),
			8884 => std_logic_vector(to_unsigned(40, 8)),
			8885 => std_logic_vector(to_unsigned(147, 8)),
			8886 => std_logic_vector(to_unsigned(231, 8)),
			8887 => std_logic_vector(to_unsigned(190, 8)),
			8888 => std_logic_vector(to_unsigned(142, 8)),
			8889 => std_logic_vector(to_unsigned(187, 8)),
			8890 => std_logic_vector(to_unsigned(12, 8)),
			8891 => std_logic_vector(to_unsigned(177, 8)),
			8892 => std_logic_vector(to_unsigned(88, 8)),
			8893 => std_logic_vector(to_unsigned(225, 8)),
			8894 => std_logic_vector(to_unsigned(90, 8)),
			8895 => std_logic_vector(to_unsigned(174, 8)),
			8896 => std_logic_vector(to_unsigned(42, 8)),
			8897 => std_logic_vector(to_unsigned(93, 8)),
			8898 => std_logic_vector(to_unsigned(26, 8)),
			8899 => std_logic_vector(to_unsigned(233, 8)),
			8900 => std_logic_vector(to_unsigned(37, 8)),
			8901 => std_logic_vector(to_unsigned(13, 8)),
			8902 => std_logic_vector(to_unsigned(242, 8)),
			8903 => std_logic_vector(to_unsigned(224, 8)),
			8904 => std_logic_vector(to_unsigned(112, 8)),
			8905 => std_logic_vector(to_unsigned(13, 8)),
			8906 => std_logic_vector(to_unsigned(245, 8)),
			8907 => std_logic_vector(to_unsigned(198, 8)),
			8908 => std_logic_vector(to_unsigned(14, 8)),
			8909 => std_logic_vector(to_unsigned(48, 8)),
			8910 => std_logic_vector(to_unsigned(243, 8)),
			8911 => std_logic_vector(to_unsigned(18, 8)),
			8912 => std_logic_vector(to_unsigned(84, 8)),
			8913 => std_logic_vector(to_unsigned(250, 8)),
			8914 => std_logic_vector(to_unsigned(85, 8)),
			8915 => std_logic_vector(to_unsigned(135, 8)),
			8916 => std_logic_vector(to_unsigned(57, 8)),
			8917 => std_logic_vector(to_unsigned(208, 8)),
			8918 => std_logic_vector(to_unsigned(28, 8)),
			8919 => std_logic_vector(to_unsigned(134, 8)),
			8920 => std_logic_vector(to_unsigned(174, 8)),
			8921 => std_logic_vector(to_unsigned(182, 8)),
			8922 => std_logic_vector(to_unsigned(244, 8)),
			8923 => std_logic_vector(to_unsigned(202, 8)),
			8924 => std_logic_vector(to_unsigned(141, 8)),
			8925 => std_logic_vector(to_unsigned(198, 8)),
			8926 => std_logic_vector(to_unsigned(103, 8)),
			8927 => std_logic_vector(to_unsigned(15, 8)),
			8928 => std_logic_vector(to_unsigned(39, 8)),
			8929 => std_logic_vector(to_unsigned(49, 8)),
			8930 => std_logic_vector(to_unsigned(21, 8)),
			8931 => std_logic_vector(to_unsigned(133, 8)),
			8932 => std_logic_vector(to_unsigned(185, 8)),
			8933 => std_logic_vector(to_unsigned(232, 8)),
			8934 => std_logic_vector(to_unsigned(34, 8)),
			8935 => std_logic_vector(to_unsigned(234, 8)),
			8936 => std_logic_vector(to_unsigned(227, 8)),
			8937 => std_logic_vector(to_unsigned(61, 8)),
			8938 => std_logic_vector(to_unsigned(10, 8)),
			8939 => std_logic_vector(to_unsigned(154, 8)),
			8940 => std_logic_vector(to_unsigned(139, 8)),
			8941 => std_logic_vector(to_unsigned(68, 8)),
			8942 => std_logic_vector(to_unsigned(232, 8)),
			8943 => std_logic_vector(to_unsigned(234, 8)),
			8944 => std_logic_vector(to_unsigned(1, 8)),
			8945 => std_logic_vector(to_unsigned(128, 8)),
			8946 => std_logic_vector(to_unsigned(103, 8)),
			8947 => std_logic_vector(to_unsigned(21, 8)),
			8948 => std_logic_vector(to_unsigned(40, 8)),
			8949 => std_logic_vector(to_unsigned(217, 8)),
			8950 => std_logic_vector(to_unsigned(4, 8)),
			8951 => std_logic_vector(to_unsigned(168, 8)),
			8952 => std_logic_vector(to_unsigned(143, 8)),
			8953 => std_logic_vector(to_unsigned(153, 8)),
			8954 => std_logic_vector(to_unsigned(161, 8)),
			8955 => std_logic_vector(to_unsigned(255, 8)),
			8956 => std_logic_vector(to_unsigned(186, 8)),
			8957 => std_logic_vector(to_unsigned(220, 8)),
			8958 => std_logic_vector(to_unsigned(183, 8)),
			8959 => std_logic_vector(to_unsigned(157, 8)),
			8960 => std_logic_vector(to_unsigned(211, 8)),
			8961 => std_logic_vector(to_unsigned(7, 8)),
			8962 => std_logic_vector(to_unsigned(243, 8)),
			8963 => std_logic_vector(to_unsigned(135, 8)),
			8964 => std_logic_vector(to_unsigned(152, 8)),
			8965 => std_logic_vector(to_unsigned(193, 8)),
			8966 => std_logic_vector(to_unsigned(221, 8)),
			8967 => std_logic_vector(to_unsigned(185, 8)),
			8968 => std_logic_vector(to_unsigned(177, 8)),
			8969 => std_logic_vector(to_unsigned(221, 8)),
			8970 => std_logic_vector(to_unsigned(237, 8)),
			8971 => std_logic_vector(to_unsigned(253, 8)),
			8972 => std_logic_vector(to_unsigned(76, 8)),
			8973 => std_logic_vector(to_unsigned(204, 8)),
			8974 => std_logic_vector(to_unsigned(216, 8)),
			8975 => std_logic_vector(to_unsigned(208, 8)),
			8976 => std_logic_vector(to_unsigned(68, 8)),
			8977 => std_logic_vector(to_unsigned(76, 8)),
			8978 => std_logic_vector(to_unsigned(39, 8)),
			8979 => std_logic_vector(to_unsigned(119, 8)),
			8980 => std_logic_vector(to_unsigned(125, 8)),
			8981 => std_logic_vector(to_unsigned(90, 8)),
			8982 => std_logic_vector(to_unsigned(133, 8)),
			8983 => std_logic_vector(to_unsigned(67, 8)),
			8984 => std_logic_vector(to_unsigned(237, 8)),
			8985 => std_logic_vector(to_unsigned(135, 8)),
			8986 => std_logic_vector(to_unsigned(199, 8)),
			8987 => std_logic_vector(to_unsigned(112, 8)),
			8988 => std_logic_vector(to_unsigned(65, 8)),
			8989 => std_logic_vector(to_unsigned(115, 8)),
			8990 => std_logic_vector(to_unsigned(200, 8)),
			8991 => std_logic_vector(to_unsigned(52, 8)),
			8992 => std_logic_vector(to_unsigned(162, 8)),
			8993 => std_logic_vector(to_unsigned(96, 8)),
			8994 => std_logic_vector(to_unsigned(39, 8)),
			8995 => std_logic_vector(to_unsigned(222, 8)),
			8996 => std_logic_vector(to_unsigned(195, 8)),
			8997 => std_logic_vector(to_unsigned(58, 8)),
			8998 => std_logic_vector(to_unsigned(15, 8)),
			8999 => std_logic_vector(to_unsigned(86, 8)),
			9000 => std_logic_vector(to_unsigned(142, 8)),
			9001 => std_logic_vector(to_unsigned(188, 8)),
			9002 => std_logic_vector(to_unsigned(129, 8)),
			9003 => std_logic_vector(to_unsigned(45, 8)),
			9004 => std_logic_vector(to_unsigned(152, 8)),
			9005 => std_logic_vector(to_unsigned(11, 8)),
			9006 => std_logic_vector(to_unsigned(76, 8)),
			9007 => std_logic_vector(to_unsigned(94, 8)),
			9008 => std_logic_vector(to_unsigned(66, 8)),
			9009 => std_logic_vector(to_unsigned(25, 8)),
			9010 => std_logic_vector(to_unsigned(100, 8)),
			9011 => std_logic_vector(to_unsigned(167, 8)),
			9012 => std_logic_vector(to_unsigned(165, 8)),
			9013 => std_logic_vector(to_unsigned(24, 8)),
			9014 => std_logic_vector(to_unsigned(58, 8)),
			9015 => std_logic_vector(to_unsigned(125, 8)),
			9016 => std_logic_vector(to_unsigned(157, 8)),
			9017 => std_logic_vector(to_unsigned(71, 8)),
			9018 => std_logic_vector(to_unsigned(165, 8)),
			9019 => std_logic_vector(to_unsigned(5, 8)),
			9020 => std_logic_vector(to_unsigned(187, 8)),
			9021 => std_logic_vector(to_unsigned(238, 8)),
			9022 => std_logic_vector(to_unsigned(82, 8)),
			9023 => std_logic_vector(to_unsigned(99, 8)),
			9024 => std_logic_vector(to_unsigned(114, 8)),
			9025 => std_logic_vector(to_unsigned(170, 8)),
			9026 => std_logic_vector(to_unsigned(142, 8)),
			9027 => std_logic_vector(to_unsigned(236, 8)),
			9028 => std_logic_vector(to_unsigned(19, 8)),
			9029 => std_logic_vector(to_unsigned(221, 8)),
			9030 => std_logic_vector(to_unsigned(56, 8)),
			9031 => std_logic_vector(to_unsigned(45, 8)),
			9032 => std_logic_vector(to_unsigned(22, 8)),
			9033 => std_logic_vector(to_unsigned(180, 8)),
			9034 => std_logic_vector(to_unsigned(12, 8)),
			9035 => std_logic_vector(to_unsigned(46, 8)),
			9036 => std_logic_vector(to_unsigned(13, 8)),
			9037 => std_logic_vector(to_unsigned(227, 8)),
			9038 => std_logic_vector(to_unsigned(201, 8)),
			9039 => std_logic_vector(to_unsigned(148, 8)),
			9040 => std_logic_vector(to_unsigned(34, 8)),
			9041 => std_logic_vector(to_unsigned(178, 8)),
			9042 => std_logic_vector(to_unsigned(202, 8)),
			9043 => std_logic_vector(to_unsigned(24, 8)),
			9044 => std_logic_vector(to_unsigned(80, 8)),
			9045 => std_logic_vector(to_unsigned(45, 8)),
			9046 => std_logic_vector(to_unsigned(52, 8)),
			9047 => std_logic_vector(to_unsigned(210, 8)),
			9048 => std_logic_vector(to_unsigned(17, 8)),
			9049 => std_logic_vector(to_unsigned(193, 8)),
			9050 => std_logic_vector(to_unsigned(86, 8)),
			9051 => std_logic_vector(to_unsigned(121, 8)),
			9052 => std_logic_vector(to_unsigned(225, 8)),
			9053 => std_logic_vector(to_unsigned(26, 8)),
			9054 => std_logic_vector(to_unsigned(228, 8)),
			9055 => std_logic_vector(to_unsigned(123, 8)),
			9056 => std_logic_vector(to_unsigned(221, 8)),
			9057 => std_logic_vector(to_unsigned(221, 8)),
			9058 => std_logic_vector(to_unsigned(81, 8)),
			9059 => std_logic_vector(to_unsigned(225, 8)),
			9060 => std_logic_vector(to_unsigned(235, 8)),
			9061 => std_logic_vector(to_unsigned(199, 8)),
			9062 => std_logic_vector(to_unsigned(194, 8)),
			9063 => std_logic_vector(to_unsigned(35, 8)),
			9064 => std_logic_vector(to_unsigned(37, 8)),
			9065 => std_logic_vector(to_unsigned(85, 8)),
			9066 => std_logic_vector(to_unsigned(72, 8)),
			9067 => std_logic_vector(to_unsigned(47, 8)),
			9068 => std_logic_vector(to_unsigned(70, 8)),
			9069 => std_logic_vector(to_unsigned(45, 8)),
			9070 => std_logic_vector(to_unsigned(124, 8)),
			9071 => std_logic_vector(to_unsigned(199, 8)),
			9072 => std_logic_vector(to_unsigned(49, 8)),
			9073 => std_logic_vector(to_unsigned(156, 8)),
			9074 => std_logic_vector(to_unsigned(225, 8)),
			9075 => std_logic_vector(to_unsigned(191, 8)),
			9076 => std_logic_vector(to_unsigned(60, 8)),
			9077 => std_logic_vector(to_unsigned(216, 8)),
			9078 => std_logic_vector(to_unsigned(31, 8)),
			9079 => std_logic_vector(to_unsigned(56, 8)),
			9080 => std_logic_vector(to_unsigned(34, 8)),
			9081 => std_logic_vector(to_unsigned(49, 8)),
			9082 => std_logic_vector(to_unsigned(194, 8)),
			9083 => std_logic_vector(to_unsigned(196, 8)),
			9084 => std_logic_vector(to_unsigned(254, 8)),
			9085 => std_logic_vector(to_unsigned(133, 8)),
			9086 => std_logic_vector(to_unsigned(247, 8)),
			9087 => std_logic_vector(to_unsigned(163, 8)),
			9088 => std_logic_vector(to_unsigned(250, 8)),
			9089 => std_logic_vector(to_unsigned(177, 8)),
			9090 => std_logic_vector(to_unsigned(123, 8)),
			9091 => std_logic_vector(to_unsigned(227, 8)),
			9092 => std_logic_vector(to_unsigned(95, 8)),
			9093 => std_logic_vector(to_unsigned(236, 8)),
			9094 => std_logic_vector(to_unsigned(42, 8)),
			9095 => std_logic_vector(to_unsigned(208, 8)),
			9096 => std_logic_vector(to_unsigned(155, 8)),
			9097 => std_logic_vector(to_unsigned(156, 8)),
			9098 => std_logic_vector(to_unsigned(224, 8)),
			9099 => std_logic_vector(to_unsigned(82, 8)),
			9100 => std_logic_vector(to_unsigned(207, 8)),
			9101 => std_logic_vector(to_unsigned(223, 8)),
			9102 => std_logic_vector(to_unsigned(251, 8)),
			9103 => std_logic_vector(to_unsigned(76, 8)),
			9104 => std_logic_vector(to_unsigned(186, 8)),
			9105 => std_logic_vector(to_unsigned(130, 8)),
			9106 => std_logic_vector(to_unsigned(63, 8)),
			9107 => std_logic_vector(to_unsigned(150, 8)),
			9108 => std_logic_vector(to_unsigned(211, 8)),
			9109 => std_logic_vector(to_unsigned(200, 8)),
			9110 => std_logic_vector(to_unsigned(178, 8)),
			9111 => std_logic_vector(to_unsigned(217, 8)),
			9112 => std_logic_vector(to_unsigned(42, 8)),
			9113 => std_logic_vector(to_unsigned(174, 8)),
			9114 => std_logic_vector(to_unsigned(22, 8)),
			9115 => std_logic_vector(to_unsigned(28, 8)),
			9116 => std_logic_vector(to_unsigned(32, 8)),
			9117 => std_logic_vector(to_unsigned(214, 8)),
			9118 => std_logic_vector(to_unsigned(109, 8)),
			9119 => std_logic_vector(to_unsigned(45, 8)),
			9120 => std_logic_vector(to_unsigned(247, 8)),
			9121 => std_logic_vector(to_unsigned(86, 8)),
			9122 => std_logic_vector(to_unsigned(92, 8)),
			9123 => std_logic_vector(to_unsigned(58, 8)),
			9124 => std_logic_vector(to_unsigned(10, 8)),
			9125 => std_logic_vector(to_unsigned(184, 8)),
			9126 => std_logic_vector(to_unsigned(5, 8)),
			9127 => std_logic_vector(to_unsigned(167, 8)),
			9128 => std_logic_vector(to_unsigned(230, 8)),
			9129 => std_logic_vector(to_unsigned(204, 8)),
			9130 => std_logic_vector(to_unsigned(39, 8)),
			9131 => std_logic_vector(to_unsigned(174, 8)),
			9132 => std_logic_vector(to_unsigned(105, 8)),
			9133 => std_logic_vector(to_unsigned(73, 8)),
			9134 => std_logic_vector(to_unsigned(20, 8)),
			9135 => std_logic_vector(to_unsigned(130, 8)),
			9136 => std_logic_vector(to_unsigned(119, 8)),
			9137 => std_logic_vector(to_unsigned(100, 8)),
			9138 => std_logic_vector(to_unsigned(60, 8)),
			9139 => std_logic_vector(to_unsigned(251, 8)),
			9140 => std_logic_vector(to_unsigned(244, 8)),
			9141 => std_logic_vector(to_unsigned(149, 8)),
			9142 => std_logic_vector(to_unsigned(41, 8)),
			9143 => std_logic_vector(to_unsigned(79, 8)),
			9144 => std_logic_vector(to_unsigned(83, 8)),
			9145 => std_logic_vector(to_unsigned(242, 8)),
			9146 => std_logic_vector(to_unsigned(249, 8)),
			9147 => std_logic_vector(to_unsigned(232, 8)),
			9148 => std_logic_vector(to_unsigned(164, 8)),
			9149 => std_logic_vector(to_unsigned(146, 8)),
			9150 => std_logic_vector(to_unsigned(180, 8)),
			9151 => std_logic_vector(to_unsigned(117, 8)),
			9152 => std_logic_vector(to_unsigned(13, 8)),
			9153 => std_logic_vector(to_unsigned(241, 8)),
			9154 => std_logic_vector(to_unsigned(230, 8)),
			9155 => std_logic_vector(to_unsigned(215, 8)),
			9156 => std_logic_vector(to_unsigned(205, 8)),
			9157 => std_logic_vector(to_unsigned(120, 8)),
			9158 => std_logic_vector(to_unsigned(78, 8)),
			9159 => std_logic_vector(to_unsigned(166, 8)),
			9160 => std_logic_vector(to_unsigned(128, 8)),
			9161 => std_logic_vector(to_unsigned(144, 8)),
			9162 => std_logic_vector(to_unsigned(136, 8)),
			9163 => std_logic_vector(to_unsigned(143, 8)),
			9164 => std_logic_vector(to_unsigned(23, 8)),
			9165 => std_logic_vector(to_unsigned(181, 8)),
			9166 => std_logic_vector(to_unsigned(100, 8)),
			9167 => std_logic_vector(to_unsigned(63, 8)),
			9168 => std_logic_vector(to_unsigned(46, 8)),
			9169 => std_logic_vector(to_unsigned(203, 8)),
			9170 => std_logic_vector(to_unsigned(92, 8)),
			9171 => std_logic_vector(to_unsigned(25, 8)),
			9172 => std_logic_vector(to_unsigned(185, 8)),
			9173 => std_logic_vector(to_unsigned(223, 8)),
			9174 => std_logic_vector(to_unsigned(132, 8)),
			9175 => std_logic_vector(to_unsigned(151, 8)),
			9176 => std_logic_vector(to_unsigned(22, 8)),
			9177 => std_logic_vector(to_unsigned(251, 8)),
			9178 => std_logic_vector(to_unsigned(124, 8)),
			9179 => std_logic_vector(to_unsigned(244, 8)),
			9180 => std_logic_vector(to_unsigned(12, 8)),
			9181 => std_logic_vector(to_unsigned(7, 8)),
			9182 => std_logic_vector(to_unsigned(51, 8)),
			9183 => std_logic_vector(to_unsigned(191, 8)),
			9184 => std_logic_vector(to_unsigned(42, 8)),
			9185 => std_logic_vector(to_unsigned(109, 8)),
			9186 => std_logic_vector(to_unsigned(35, 8)),
			9187 => std_logic_vector(to_unsigned(75, 8)),
			9188 => std_logic_vector(to_unsigned(185, 8)),
			9189 => std_logic_vector(to_unsigned(33, 8)),
			9190 => std_logic_vector(to_unsigned(38, 8)),
			9191 => std_logic_vector(to_unsigned(67, 8)),
			9192 => std_logic_vector(to_unsigned(150, 8)),
			9193 => std_logic_vector(to_unsigned(108, 8)),
			9194 => std_logic_vector(to_unsigned(179, 8)),
			9195 => std_logic_vector(to_unsigned(189, 8)),
			9196 => std_logic_vector(to_unsigned(15, 8)),
			9197 => std_logic_vector(to_unsigned(35, 8)),
			9198 => std_logic_vector(to_unsigned(75, 8)),
			9199 => std_logic_vector(to_unsigned(73, 8)),
			9200 => std_logic_vector(to_unsigned(160, 8)),
			9201 => std_logic_vector(to_unsigned(218, 8)),
			9202 => std_logic_vector(to_unsigned(220, 8)),
			9203 => std_logic_vector(to_unsigned(89, 8)),
			9204 => std_logic_vector(to_unsigned(145, 8)),
			9205 => std_logic_vector(to_unsigned(51, 8)),
			9206 => std_logic_vector(to_unsigned(96, 8)),
			9207 => std_logic_vector(to_unsigned(248, 8)),
			9208 => std_logic_vector(to_unsigned(159, 8)),
			9209 => std_logic_vector(to_unsigned(124, 8)),
			9210 => std_logic_vector(to_unsigned(11, 8)),
			9211 => std_logic_vector(to_unsigned(96, 8)),
			9212 => std_logic_vector(to_unsigned(251, 8)),
			9213 => std_logic_vector(to_unsigned(96, 8)),
			9214 => std_logic_vector(to_unsigned(17, 8)),
			9215 => std_logic_vector(to_unsigned(228, 8)),
			9216 => std_logic_vector(to_unsigned(219, 8)),
			9217 => std_logic_vector(to_unsigned(18, 8)),
			9218 => std_logic_vector(to_unsigned(185, 8)),
			9219 => std_logic_vector(to_unsigned(137, 8)),
			9220 => std_logic_vector(to_unsigned(192, 8)),
			9221 => std_logic_vector(to_unsigned(110, 8)),
			9222 => std_logic_vector(to_unsigned(197, 8)),
			9223 => std_logic_vector(to_unsigned(1, 8)),
			9224 => std_logic_vector(to_unsigned(34, 8)),
			9225 => std_logic_vector(to_unsigned(179, 8)),
			9226 => std_logic_vector(to_unsigned(240, 8)),
			9227 => std_logic_vector(to_unsigned(116, 8)),
			9228 => std_logic_vector(to_unsigned(209, 8)),
			9229 => std_logic_vector(to_unsigned(194, 8)),
			9230 => std_logic_vector(to_unsigned(198, 8)),
			9231 => std_logic_vector(to_unsigned(33, 8)),
			9232 => std_logic_vector(to_unsigned(92, 8)),
			9233 => std_logic_vector(to_unsigned(229, 8)),
			9234 => std_logic_vector(to_unsigned(51, 8)),
			9235 => std_logic_vector(to_unsigned(155, 8)),
			9236 => std_logic_vector(to_unsigned(42, 8)),
			9237 => std_logic_vector(to_unsigned(136, 8)),
			9238 => std_logic_vector(to_unsigned(66, 8)),
			9239 => std_logic_vector(to_unsigned(243, 8)),
			9240 => std_logic_vector(to_unsigned(33, 8)),
			9241 => std_logic_vector(to_unsigned(232, 8)),
			9242 => std_logic_vector(to_unsigned(14, 8)),
			9243 => std_logic_vector(to_unsigned(50, 8)),
			9244 => std_logic_vector(to_unsigned(110, 8)),
			9245 => std_logic_vector(to_unsigned(214, 8)),
			9246 => std_logic_vector(to_unsigned(148, 8)),
			9247 => std_logic_vector(to_unsigned(109, 8)),
			9248 => std_logic_vector(to_unsigned(98, 8)),
			9249 => std_logic_vector(to_unsigned(72, 8)),
			9250 => std_logic_vector(to_unsigned(83, 8)),
			9251 => std_logic_vector(to_unsigned(45, 8)),
			9252 => std_logic_vector(to_unsigned(51, 8)),
			9253 => std_logic_vector(to_unsigned(188, 8)),
			9254 => std_logic_vector(to_unsigned(177, 8)),
			9255 => std_logic_vector(to_unsigned(154, 8)),
			9256 => std_logic_vector(to_unsigned(123, 8)),
			9257 => std_logic_vector(to_unsigned(226, 8)),
			9258 => std_logic_vector(to_unsigned(210, 8)),
			9259 => std_logic_vector(to_unsigned(54, 8)),
			9260 => std_logic_vector(to_unsigned(33, 8)),
			9261 => std_logic_vector(to_unsigned(144, 8)),
			9262 => std_logic_vector(to_unsigned(254, 8)),
			9263 => std_logic_vector(to_unsigned(120, 8)),
			9264 => std_logic_vector(to_unsigned(33, 8)),
			9265 => std_logic_vector(to_unsigned(218, 8)),
			9266 => std_logic_vector(to_unsigned(80, 8)),
			9267 => std_logic_vector(to_unsigned(7, 8)),
			9268 => std_logic_vector(to_unsigned(61, 8)),
			9269 => std_logic_vector(to_unsigned(119, 8)),
			9270 => std_logic_vector(to_unsigned(48, 8)),
			9271 => std_logic_vector(to_unsigned(151, 8)),
			9272 => std_logic_vector(to_unsigned(250, 8)),
			9273 => std_logic_vector(to_unsigned(210, 8)),
			9274 => std_logic_vector(to_unsigned(178, 8)),
			9275 => std_logic_vector(to_unsigned(199, 8)),
			9276 => std_logic_vector(to_unsigned(32, 8)),
			9277 => std_logic_vector(to_unsigned(71, 8)),
			9278 => std_logic_vector(to_unsigned(186, 8)),
			9279 => std_logic_vector(to_unsigned(83, 8)),
			9280 => std_logic_vector(to_unsigned(226, 8)),
			9281 => std_logic_vector(to_unsigned(60, 8)),
			9282 => std_logic_vector(to_unsigned(155, 8)),
			9283 => std_logic_vector(to_unsigned(204, 8)),
			9284 => std_logic_vector(to_unsigned(196, 8)),
			9285 => std_logic_vector(to_unsigned(227, 8)),
			9286 => std_logic_vector(to_unsigned(240, 8)),
			9287 => std_logic_vector(to_unsigned(249, 8)),
			9288 => std_logic_vector(to_unsigned(228, 8)),
			9289 => std_logic_vector(to_unsigned(161, 8)),
			9290 => std_logic_vector(to_unsigned(93, 8)),
			9291 => std_logic_vector(to_unsigned(114, 8)),
			9292 => std_logic_vector(to_unsigned(198, 8)),
			9293 => std_logic_vector(to_unsigned(85, 8)),
			9294 => std_logic_vector(to_unsigned(88, 8)),
			9295 => std_logic_vector(to_unsigned(29, 8)),
			9296 => std_logic_vector(to_unsigned(128, 8)),
			9297 => std_logic_vector(to_unsigned(160, 8)),
			9298 => std_logic_vector(to_unsigned(220, 8)),
			9299 => std_logic_vector(to_unsigned(191, 8)),
			9300 => std_logic_vector(to_unsigned(196, 8)),
			9301 => std_logic_vector(to_unsigned(51, 8)),
			9302 => std_logic_vector(to_unsigned(229, 8)),
			9303 => std_logic_vector(to_unsigned(82, 8)),
			9304 => std_logic_vector(to_unsigned(114, 8)),
			9305 => std_logic_vector(to_unsigned(231, 8)),
			9306 => std_logic_vector(to_unsigned(80, 8)),
			9307 => std_logic_vector(to_unsigned(34, 8)),
			9308 => std_logic_vector(to_unsigned(80, 8)),
			9309 => std_logic_vector(to_unsigned(199, 8)),
			9310 => std_logic_vector(to_unsigned(240, 8)),
			9311 => std_logic_vector(to_unsigned(246, 8)),
			9312 => std_logic_vector(to_unsigned(184, 8)),
			9313 => std_logic_vector(to_unsigned(89, 8)),
			9314 => std_logic_vector(to_unsigned(66, 8)),
			9315 => std_logic_vector(to_unsigned(211, 8)),
			9316 => std_logic_vector(to_unsigned(148, 8)),
			9317 => std_logic_vector(to_unsigned(99, 8)),
			9318 => std_logic_vector(to_unsigned(149, 8)),
			9319 => std_logic_vector(to_unsigned(79, 8)),
			9320 => std_logic_vector(to_unsigned(124, 8)),
			9321 => std_logic_vector(to_unsigned(15, 8)),
			9322 => std_logic_vector(to_unsigned(230, 8)),
			9323 => std_logic_vector(to_unsigned(105, 8)),
			9324 => std_logic_vector(to_unsigned(213, 8)),
			9325 => std_logic_vector(to_unsigned(216, 8)),
			9326 => std_logic_vector(to_unsigned(215, 8)),
			9327 => std_logic_vector(to_unsigned(47, 8)),
			9328 => std_logic_vector(to_unsigned(208, 8)),
			9329 => std_logic_vector(to_unsigned(26, 8)),
			9330 => std_logic_vector(to_unsigned(211, 8)),
			9331 => std_logic_vector(to_unsigned(38, 8)),
			9332 => std_logic_vector(to_unsigned(172, 8)),
			9333 => std_logic_vector(to_unsigned(36, 8)),
			9334 => std_logic_vector(to_unsigned(127, 8)),
			9335 => std_logic_vector(to_unsigned(37, 8)),
			9336 => std_logic_vector(to_unsigned(142, 8)),
			9337 => std_logic_vector(to_unsigned(194, 8)),
			9338 => std_logic_vector(to_unsigned(171, 8)),
			9339 => std_logic_vector(to_unsigned(45, 8)),
			9340 => std_logic_vector(to_unsigned(117, 8)),
			9341 => std_logic_vector(to_unsigned(16, 8)),
			9342 => std_logic_vector(to_unsigned(133, 8)),
			9343 => std_logic_vector(to_unsigned(165, 8)),
			9344 => std_logic_vector(to_unsigned(143, 8)),
			9345 => std_logic_vector(to_unsigned(12, 8)),
			9346 => std_logic_vector(to_unsigned(86, 8)),
			9347 => std_logic_vector(to_unsigned(209, 8)),
			9348 => std_logic_vector(to_unsigned(208, 8)),
			9349 => std_logic_vector(to_unsigned(124, 8)),
			9350 => std_logic_vector(to_unsigned(175, 8)),
			9351 => std_logic_vector(to_unsigned(132, 8)),
			9352 => std_logic_vector(to_unsigned(88, 8)),
			9353 => std_logic_vector(to_unsigned(183, 8)),
			9354 => std_logic_vector(to_unsigned(94, 8)),
			9355 => std_logic_vector(to_unsigned(44, 8)),
			9356 => std_logic_vector(to_unsigned(93, 8)),
			9357 => std_logic_vector(to_unsigned(35, 8)),
			9358 => std_logic_vector(to_unsigned(113, 8)),
			9359 => std_logic_vector(to_unsigned(234, 8)),
			9360 => std_logic_vector(to_unsigned(63, 8)),
			9361 => std_logic_vector(to_unsigned(153, 8)),
			9362 => std_logic_vector(to_unsigned(0, 8)),
			9363 => std_logic_vector(to_unsigned(171, 8)),
			9364 => std_logic_vector(to_unsigned(226, 8)),
			9365 => std_logic_vector(to_unsigned(211, 8)),
			9366 => std_logic_vector(to_unsigned(147, 8)),
			9367 => std_logic_vector(to_unsigned(176, 8)),
			9368 => std_logic_vector(to_unsigned(59, 8)),
			9369 => std_logic_vector(to_unsigned(60, 8)),
			9370 => std_logic_vector(to_unsigned(40, 8)),
			9371 => std_logic_vector(to_unsigned(41, 8)),
			9372 => std_logic_vector(to_unsigned(65, 8)),
			9373 => std_logic_vector(to_unsigned(63, 8)),
			9374 => std_logic_vector(to_unsigned(119, 8)),
			9375 => std_logic_vector(to_unsigned(74, 8)),
			9376 => std_logic_vector(to_unsigned(201, 8)),
			9377 => std_logic_vector(to_unsigned(44, 8)),
			9378 => std_logic_vector(to_unsigned(136, 8)),
			9379 => std_logic_vector(to_unsigned(118, 8)),
			9380 => std_logic_vector(to_unsigned(138, 8)),
			9381 => std_logic_vector(to_unsigned(239, 8)),
			9382 => std_logic_vector(to_unsigned(57, 8)),
			9383 => std_logic_vector(to_unsigned(244, 8)),
			9384 => std_logic_vector(to_unsigned(40, 8)),
			9385 => std_logic_vector(to_unsigned(31, 8)),
			9386 => std_logic_vector(to_unsigned(39, 8)),
			9387 => std_logic_vector(to_unsigned(81, 8)),
			9388 => std_logic_vector(to_unsigned(172, 8)),
			9389 => std_logic_vector(to_unsigned(177, 8)),
			9390 => std_logic_vector(to_unsigned(190, 8)),
			9391 => std_logic_vector(to_unsigned(44, 8)),
			9392 => std_logic_vector(to_unsigned(164, 8)),
			9393 => std_logic_vector(to_unsigned(49, 8)),
			9394 => std_logic_vector(to_unsigned(35, 8)),
			9395 => std_logic_vector(to_unsigned(115, 8)),
			9396 => std_logic_vector(to_unsigned(236, 8)),
			9397 => std_logic_vector(to_unsigned(138, 8)),
			9398 => std_logic_vector(to_unsigned(100, 8)),
			9399 => std_logic_vector(to_unsigned(118, 8)),
			9400 => std_logic_vector(to_unsigned(210, 8)),
			9401 => std_logic_vector(to_unsigned(147, 8)),
			9402 => std_logic_vector(to_unsigned(78, 8)),
			9403 => std_logic_vector(to_unsigned(33, 8)),
			9404 => std_logic_vector(to_unsigned(112, 8)),
			9405 => std_logic_vector(to_unsigned(248, 8)),
			9406 => std_logic_vector(to_unsigned(7, 8)),
			9407 => std_logic_vector(to_unsigned(136, 8)),
			9408 => std_logic_vector(to_unsigned(139, 8)),
			9409 => std_logic_vector(to_unsigned(158, 8)),
			9410 => std_logic_vector(to_unsigned(33, 8)),
			9411 => std_logic_vector(to_unsigned(149, 8)),
			9412 => std_logic_vector(to_unsigned(6, 8)),
			9413 => std_logic_vector(to_unsigned(137, 8)),
			9414 => std_logic_vector(to_unsigned(68, 8)),
			9415 => std_logic_vector(to_unsigned(165, 8)),
			9416 => std_logic_vector(to_unsigned(3, 8)),
			9417 => std_logic_vector(to_unsigned(90, 8)),
			9418 => std_logic_vector(to_unsigned(187, 8)),
			9419 => std_logic_vector(to_unsigned(198, 8)),
			9420 => std_logic_vector(to_unsigned(178, 8)),
			9421 => std_logic_vector(to_unsigned(81, 8)),
			9422 => std_logic_vector(to_unsigned(138, 8)),
			9423 => std_logic_vector(to_unsigned(90, 8)),
			9424 => std_logic_vector(to_unsigned(229, 8)),
			9425 => std_logic_vector(to_unsigned(58, 8)),
			9426 => std_logic_vector(to_unsigned(38, 8)),
			9427 => std_logic_vector(to_unsigned(82, 8)),
			9428 => std_logic_vector(to_unsigned(72, 8)),
			9429 => std_logic_vector(to_unsigned(98, 8)),
			9430 => std_logic_vector(to_unsigned(111, 8)),
			9431 => std_logic_vector(to_unsigned(104, 8)),
			9432 => std_logic_vector(to_unsigned(62, 8)),
			9433 => std_logic_vector(to_unsigned(240, 8)),
			9434 => std_logic_vector(to_unsigned(75, 8)),
			9435 => std_logic_vector(to_unsigned(181, 8)),
			9436 => std_logic_vector(to_unsigned(35, 8)),
			9437 => std_logic_vector(to_unsigned(53, 8)),
			9438 => std_logic_vector(to_unsigned(43, 8)),
			9439 => std_logic_vector(to_unsigned(124, 8)),
			9440 => std_logic_vector(to_unsigned(45, 8)),
			9441 => std_logic_vector(to_unsigned(155, 8)),
			9442 => std_logic_vector(to_unsigned(8, 8)),
			9443 => std_logic_vector(to_unsigned(79, 8)),
			9444 => std_logic_vector(to_unsigned(38, 8)),
			9445 => std_logic_vector(to_unsigned(78, 8)),
			9446 => std_logic_vector(to_unsigned(243, 8)),
			9447 => std_logic_vector(to_unsigned(246, 8)),
			9448 => std_logic_vector(to_unsigned(127, 8)),
			9449 => std_logic_vector(to_unsigned(78, 8)),
			9450 => std_logic_vector(to_unsigned(174, 8)),
			9451 => std_logic_vector(to_unsigned(112, 8)),
			9452 => std_logic_vector(to_unsigned(231, 8)),
			9453 => std_logic_vector(to_unsigned(194, 8)),
			9454 => std_logic_vector(to_unsigned(26, 8)),
			9455 => std_logic_vector(to_unsigned(6, 8)),
			9456 => std_logic_vector(to_unsigned(80, 8)),
			9457 => std_logic_vector(to_unsigned(4, 8)),
			9458 => std_logic_vector(to_unsigned(68, 8)),
			9459 => std_logic_vector(to_unsigned(91, 8)),
			9460 => std_logic_vector(to_unsigned(201, 8)),
			9461 => std_logic_vector(to_unsigned(221, 8)),
			9462 => std_logic_vector(to_unsigned(140, 8)),
			9463 => std_logic_vector(to_unsigned(37, 8)),
			9464 => std_logic_vector(to_unsigned(30, 8)),
			9465 => std_logic_vector(to_unsigned(110, 8)),
			9466 => std_logic_vector(to_unsigned(226, 8)),
			9467 => std_logic_vector(to_unsigned(0, 8)),
			9468 => std_logic_vector(to_unsigned(217, 8)),
			9469 => std_logic_vector(to_unsigned(127, 8)),
			9470 => std_logic_vector(to_unsigned(167, 8)),
			9471 => std_logic_vector(to_unsigned(101, 8)),
			9472 => std_logic_vector(to_unsigned(200, 8)),
			9473 => std_logic_vector(to_unsigned(82, 8)),
			9474 => std_logic_vector(to_unsigned(123, 8)),
			9475 => std_logic_vector(to_unsigned(39, 8)),
			9476 => std_logic_vector(to_unsigned(25, 8)),
			9477 => std_logic_vector(to_unsigned(16, 8)),
			9478 => std_logic_vector(to_unsigned(167, 8)),
			9479 => std_logic_vector(to_unsigned(92, 8)),
			9480 => std_logic_vector(to_unsigned(237, 8)),
			9481 => std_logic_vector(to_unsigned(213, 8)),
			9482 => std_logic_vector(to_unsigned(222, 8)),
			9483 => std_logic_vector(to_unsigned(220, 8)),
			9484 => std_logic_vector(to_unsigned(177, 8)),
			9485 => std_logic_vector(to_unsigned(55, 8)),
			9486 => std_logic_vector(to_unsigned(253, 8)),
			9487 => std_logic_vector(to_unsigned(67, 8)),
			9488 => std_logic_vector(to_unsigned(198, 8)),
			9489 => std_logic_vector(to_unsigned(197, 8)),
			9490 => std_logic_vector(to_unsigned(40, 8)),
			9491 => std_logic_vector(to_unsigned(64, 8)),
			9492 => std_logic_vector(to_unsigned(151, 8)),
			9493 => std_logic_vector(to_unsigned(6, 8)),
			9494 => std_logic_vector(to_unsigned(84, 8)),
			9495 => std_logic_vector(to_unsigned(194, 8)),
			9496 => std_logic_vector(to_unsigned(32, 8)),
			9497 => std_logic_vector(to_unsigned(67, 8)),
			9498 => std_logic_vector(to_unsigned(70, 8)),
			9499 => std_logic_vector(to_unsigned(122, 8)),
			9500 => std_logic_vector(to_unsigned(9, 8)),
			9501 => std_logic_vector(to_unsigned(62, 8)),
			9502 => std_logic_vector(to_unsigned(102, 8)),
			9503 => std_logic_vector(to_unsigned(254, 8)),
			9504 => std_logic_vector(to_unsigned(238, 8)),
			9505 => std_logic_vector(to_unsigned(221, 8)),
			9506 => std_logic_vector(to_unsigned(0, 8)),
			9507 => std_logic_vector(to_unsigned(177, 8)),
			9508 => std_logic_vector(to_unsigned(83, 8)),
			9509 => std_logic_vector(to_unsigned(51, 8)),
			9510 => std_logic_vector(to_unsigned(139, 8)),
			9511 => std_logic_vector(to_unsigned(24, 8)),
			9512 => std_logic_vector(to_unsigned(157, 8)),
			9513 => std_logic_vector(to_unsigned(40, 8)),
			9514 => std_logic_vector(to_unsigned(95, 8)),
			9515 => std_logic_vector(to_unsigned(72, 8)),
			9516 => std_logic_vector(to_unsigned(40, 8)),
			9517 => std_logic_vector(to_unsigned(30, 8)),
			9518 => std_logic_vector(to_unsigned(168, 8)),
			9519 => std_logic_vector(to_unsigned(145, 8)),
			9520 => std_logic_vector(to_unsigned(91, 8)),
			9521 => std_logic_vector(to_unsigned(26, 8)),
			9522 => std_logic_vector(to_unsigned(191, 8)),
			9523 => std_logic_vector(to_unsigned(174, 8)),
			9524 => std_logic_vector(to_unsigned(236, 8)),
			9525 => std_logic_vector(to_unsigned(132, 8)),
			9526 => std_logic_vector(to_unsigned(161, 8)),
			9527 => std_logic_vector(to_unsigned(129, 8)),
			9528 => std_logic_vector(to_unsigned(81, 8)),
			9529 => std_logic_vector(to_unsigned(107, 8)),
			9530 => std_logic_vector(to_unsigned(17, 8)),
			9531 => std_logic_vector(to_unsigned(141, 8)),
			9532 => std_logic_vector(to_unsigned(18, 8)),
			9533 => std_logic_vector(to_unsigned(61, 8)),
			9534 => std_logic_vector(to_unsigned(42, 8)),
			9535 => std_logic_vector(to_unsigned(102, 8)),
			9536 => std_logic_vector(to_unsigned(219, 8)),
			9537 => std_logic_vector(to_unsigned(162, 8)),
			9538 => std_logic_vector(to_unsigned(111, 8)),
			9539 => std_logic_vector(to_unsigned(87, 8)),
			9540 => std_logic_vector(to_unsigned(30, 8)),
			9541 => std_logic_vector(to_unsigned(96, 8)),
			9542 => std_logic_vector(to_unsigned(74, 8)),
			9543 => std_logic_vector(to_unsigned(150, 8)),
			9544 => std_logic_vector(to_unsigned(232, 8)),
			9545 => std_logic_vector(to_unsigned(2, 8)),
			9546 => std_logic_vector(to_unsigned(218, 8)),
			9547 => std_logic_vector(to_unsigned(89, 8)),
			9548 => std_logic_vector(to_unsigned(152, 8)),
			9549 => std_logic_vector(to_unsigned(171, 8)),
			9550 => std_logic_vector(to_unsigned(233, 8)),
			9551 => std_logic_vector(to_unsigned(254, 8)),
			9552 => std_logic_vector(to_unsigned(127, 8)),
			9553 => std_logic_vector(to_unsigned(245, 8)),
			9554 => std_logic_vector(to_unsigned(95, 8)),
			9555 => std_logic_vector(to_unsigned(22, 8)),
			9556 => std_logic_vector(to_unsigned(100, 8)),
			9557 => std_logic_vector(to_unsigned(113, 8)),
			9558 => std_logic_vector(to_unsigned(146, 8)),
			9559 => std_logic_vector(to_unsigned(101, 8)),
			9560 => std_logic_vector(to_unsigned(33, 8)),
			9561 => std_logic_vector(to_unsigned(142, 8)),
			9562 => std_logic_vector(to_unsigned(140, 8)),
			9563 => std_logic_vector(to_unsigned(236, 8)),
			9564 => std_logic_vector(to_unsigned(86, 8)),
			9565 => std_logic_vector(to_unsigned(29, 8)),
			9566 => std_logic_vector(to_unsigned(43, 8)),
			9567 => std_logic_vector(to_unsigned(108, 8)),
			9568 => std_logic_vector(to_unsigned(210, 8)),
			9569 => std_logic_vector(to_unsigned(243, 8)),
			9570 => std_logic_vector(to_unsigned(10, 8)),
			9571 => std_logic_vector(to_unsigned(0, 8)),
			9572 => std_logic_vector(to_unsigned(176, 8)),
			9573 => std_logic_vector(to_unsigned(40, 8)),
			9574 => std_logic_vector(to_unsigned(188, 8)),
			9575 => std_logic_vector(to_unsigned(22, 8)),
			9576 => std_logic_vector(to_unsigned(249, 8)),
			9577 => std_logic_vector(to_unsigned(188, 8)),
			9578 => std_logic_vector(to_unsigned(28, 8)),
			9579 => std_logic_vector(to_unsigned(5, 8)),
			9580 => std_logic_vector(to_unsigned(17, 8)),
			9581 => std_logic_vector(to_unsigned(228, 8)),
			9582 => std_logic_vector(to_unsigned(94, 8)),
			9583 => std_logic_vector(to_unsigned(186, 8)),
			9584 => std_logic_vector(to_unsigned(0, 8)),
			9585 => std_logic_vector(to_unsigned(171, 8)),
			9586 => std_logic_vector(to_unsigned(22, 8)),
			9587 => std_logic_vector(to_unsigned(126, 8)),
			9588 => std_logic_vector(to_unsigned(28, 8)),
			9589 => std_logic_vector(to_unsigned(52, 8)),
			9590 => std_logic_vector(to_unsigned(55, 8)),
			9591 => std_logic_vector(to_unsigned(208, 8)),
			9592 => std_logic_vector(to_unsigned(32, 8)),
			9593 => std_logic_vector(to_unsigned(6, 8)),
			9594 => std_logic_vector(to_unsigned(147, 8)),
			9595 => std_logic_vector(to_unsigned(249, 8)),
			9596 => std_logic_vector(to_unsigned(121, 8)),
			9597 => std_logic_vector(to_unsigned(204, 8)),
			9598 => std_logic_vector(to_unsigned(42, 8)),
			9599 => std_logic_vector(to_unsigned(128, 8)),
			9600 => std_logic_vector(to_unsigned(138, 8)),
			9601 => std_logic_vector(to_unsigned(66, 8)),
			9602 => std_logic_vector(to_unsigned(197, 8)),
			9603 => std_logic_vector(to_unsigned(164, 8)),
			9604 => std_logic_vector(to_unsigned(106, 8)),
			9605 => std_logic_vector(to_unsigned(98, 8)),
			9606 => std_logic_vector(to_unsigned(214, 8)),
			9607 => std_logic_vector(to_unsigned(142, 8)),
			9608 => std_logic_vector(to_unsigned(74, 8)),
			9609 => std_logic_vector(to_unsigned(234, 8)),
			9610 => std_logic_vector(to_unsigned(102, 8)),
			9611 => std_logic_vector(to_unsigned(184, 8)),
			9612 => std_logic_vector(to_unsigned(37, 8)),
			9613 => std_logic_vector(to_unsigned(174, 8)),
			9614 => std_logic_vector(to_unsigned(129, 8)),
			9615 => std_logic_vector(to_unsigned(2, 8)),
			9616 => std_logic_vector(to_unsigned(255, 8)),
			9617 => std_logic_vector(to_unsigned(223, 8)),
			9618 => std_logic_vector(to_unsigned(112, 8)),
			9619 => std_logic_vector(to_unsigned(45, 8)),
			9620 => std_logic_vector(to_unsigned(92, 8)),
			9621 => std_logic_vector(to_unsigned(150, 8)),
			9622 => std_logic_vector(to_unsigned(57, 8)),
			9623 => std_logic_vector(to_unsigned(246, 8)),
			9624 => std_logic_vector(to_unsigned(163, 8)),
			9625 => std_logic_vector(to_unsigned(50, 8)),
			9626 => std_logic_vector(to_unsigned(2, 8)),
			9627 => std_logic_vector(to_unsigned(136, 8)),
			9628 => std_logic_vector(to_unsigned(171, 8)),
			9629 => std_logic_vector(to_unsigned(42, 8)),
			9630 => std_logic_vector(to_unsigned(145, 8)),
			9631 => std_logic_vector(to_unsigned(138, 8)),
			9632 => std_logic_vector(to_unsigned(163, 8)),
			9633 => std_logic_vector(to_unsigned(210, 8)),
			9634 => std_logic_vector(to_unsigned(129, 8)),
			9635 => std_logic_vector(to_unsigned(61, 8)),
			9636 => std_logic_vector(to_unsigned(37, 8)),
			9637 => std_logic_vector(to_unsigned(193, 8)),
			9638 => std_logic_vector(to_unsigned(221, 8)),
			9639 => std_logic_vector(to_unsigned(179, 8)),
			9640 => std_logic_vector(to_unsigned(51, 8)),
			9641 => std_logic_vector(to_unsigned(76, 8)),
			9642 => std_logic_vector(to_unsigned(70, 8)),
			9643 => std_logic_vector(to_unsigned(150, 8)),
			9644 => std_logic_vector(to_unsigned(77, 8)),
			9645 => std_logic_vector(to_unsigned(219, 8)),
			9646 => std_logic_vector(to_unsigned(36, 8)),
			9647 => std_logic_vector(to_unsigned(100, 8)),
			9648 => std_logic_vector(to_unsigned(232, 8)),
			9649 => std_logic_vector(to_unsigned(109, 8)),
			9650 => std_logic_vector(to_unsigned(148, 8)),
			9651 => std_logic_vector(to_unsigned(93, 8)),
			9652 => std_logic_vector(to_unsigned(66, 8)),
			9653 => std_logic_vector(to_unsigned(21, 8)),
			9654 => std_logic_vector(to_unsigned(182, 8)),
			9655 => std_logic_vector(to_unsigned(192, 8)),
			9656 => std_logic_vector(to_unsigned(85, 8)),
			9657 => std_logic_vector(to_unsigned(164, 8)),
			9658 => std_logic_vector(to_unsigned(177, 8)),
			9659 => std_logic_vector(to_unsigned(143, 8)),
			9660 => std_logic_vector(to_unsigned(249, 8)),
			9661 => std_logic_vector(to_unsigned(241, 8)),
			9662 => std_logic_vector(to_unsigned(88, 8)),
			9663 => std_logic_vector(to_unsigned(139, 8)),
			9664 => std_logic_vector(to_unsigned(13, 8)),
			9665 => std_logic_vector(to_unsigned(75, 8)),
			9666 => std_logic_vector(to_unsigned(42, 8)),
			9667 => std_logic_vector(to_unsigned(14, 8)),
			9668 => std_logic_vector(to_unsigned(218, 8)),
			9669 => std_logic_vector(to_unsigned(193, 8)),
			9670 => std_logic_vector(to_unsigned(202, 8)),
			9671 => std_logic_vector(to_unsigned(7, 8)),
			9672 => std_logic_vector(to_unsigned(32, 8)),
			9673 => std_logic_vector(to_unsigned(79, 8)),
			9674 => std_logic_vector(to_unsigned(176, 8)),
			9675 => std_logic_vector(to_unsigned(100, 8)),
			9676 => std_logic_vector(to_unsigned(245, 8)),
			9677 => std_logic_vector(to_unsigned(118, 8)),
			9678 => std_logic_vector(to_unsigned(233, 8)),
			9679 => std_logic_vector(to_unsigned(193, 8)),
			9680 => std_logic_vector(to_unsigned(1, 8)),
			9681 => std_logic_vector(to_unsigned(245, 8)),
			9682 => std_logic_vector(to_unsigned(89, 8)),
			9683 => std_logic_vector(to_unsigned(139, 8)),
			9684 => std_logic_vector(to_unsigned(151, 8)),
			9685 => std_logic_vector(to_unsigned(98, 8)),
			9686 => std_logic_vector(to_unsigned(204, 8)),
			9687 => std_logic_vector(to_unsigned(77, 8)),
			9688 => std_logic_vector(to_unsigned(116, 8)),
			9689 => std_logic_vector(to_unsigned(184, 8)),
			9690 => std_logic_vector(to_unsigned(186, 8)),
			9691 => std_logic_vector(to_unsigned(15, 8)),
			9692 => std_logic_vector(to_unsigned(202, 8)),
			9693 => std_logic_vector(to_unsigned(2, 8)),
			9694 => std_logic_vector(to_unsigned(37, 8)),
			9695 => std_logic_vector(to_unsigned(202, 8)),
			9696 => std_logic_vector(to_unsigned(217, 8)),
			9697 => std_logic_vector(to_unsigned(111, 8)),
			9698 => std_logic_vector(to_unsigned(35, 8)),
			9699 => std_logic_vector(to_unsigned(81, 8)),
			9700 => std_logic_vector(to_unsigned(5, 8)),
			9701 => std_logic_vector(to_unsigned(41, 8)),
			9702 => std_logic_vector(to_unsigned(86, 8)),
			9703 => std_logic_vector(to_unsigned(201, 8)),
			9704 => std_logic_vector(to_unsigned(254, 8)),
			9705 => std_logic_vector(to_unsigned(236, 8)),
			9706 => std_logic_vector(to_unsigned(108, 8)),
			9707 => std_logic_vector(to_unsigned(251, 8)),
			9708 => std_logic_vector(to_unsigned(22, 8)),
			9709 => std_logic_vector(to_unsigned(186, 8)),
			9710 => std_logic_vector(to_unsigned(152, 8)),
			9711 => std_logic_vector(to_unsigned(165, 8)),
			9712 => std_logic_vector(to_unsigned(121, 8)),
			9713 => std_logic_vector(to_unsigned(25, 8)),
			9714 => std_logic_vector(to_unsigned(168, 8)),
			9715 => std_logic_vector(to_unsigned(96, 8)),
			9716 => std_logic_vector(to_unsigned(151, 8)),
			9717 => std_logic_vector(to_unsigned(96, 8)),
			9718 => std_logic_vector(to_unsigned(60, 8)),
			9719 => std_logic_vector(to_unsigned(94, 8)),
			9720 => std_logic_vector(to_unsigned(5, 8)),
			9721 => std_logic_vector(to_unsigned(90, 8)),
			9722 => std_logic_vector(to_unsigned(172, 8)),
			9723 => std_logic_vector(to_unsigned(209, 8)),
			9724 => std_logic_vector(to_unsigned(128, 8)),
			9725 => std_logic_vector(to_unsigned(205, 8)),
			9726 => std_logic_vector(to_unsigned(49, 8)),
			9727 => std_logic_vector(to_unsigned(170, 8)),
			9728 => std_logic_vector(to_unsigned(210, 8)),
			9729 => std_logic_vector(to_unsigned(225, 8)),
			9730 => std_logic_vector(to_unsigned(187, 8)),
			9731 => std_logic_vector(to_unsigned(28, 8)),
			9732 => std_logic_vector(to_unsigned(100, 8)),
			9733 => std_logic_vector(to_unsigned(61, 8)),
			9734 => std_logic_vector(to_unsigned(6, 8)),
			9735 => std_logic_vector(to_unsigned(86, 8)),
			9736 => std_logic_vector(to_unsigned(124, 8)),
			9737 => std_logic_vector(to_unsigned(56, 8)),
			9738 => std_logic_vector(to_unsigned(110, 8)),
			9739 => std_logic_vector(to_unsigned(146, 8)),
			9740 => std_logic_vector(to_unsigned(151, 8)),
			9741 => std_logic_vector(to_unsigned(239, 8)),
			9742 => std_logic_vector(to_unsigned(158, 8)),
			9743 => std_logic_vector(to_unsigned(56, 8)),
			9744 => std_logic_vector(to_unsigned(182, 8)),
			9745 => std_logic_vector(to_unsigned(83, 8)),
			9746 => std_logic_vector(to_unsigned(151, 8)),
			9747 => std_logic_vector(to_unsigned(166, 8)),
			9748 => std_logic_vector(to_unsigned(166, 8)),
			9749 => std_logic_vector(to_unsigned(43, 8)),
			9750 => std_logic_vector(to_unsigned(243, 8)),
			9751 => std_logic_vector(to_unsigned(58, 8)),
			9752 => std_logic_vector(to_unsigned(209, 8)),
			9753 => std_logic_vector(to_unsigned(11, 8)),
			9754 => std_logic_vector(to_unsigned(173, 8)),
			9755 => std_logic_vector(to_unsigned(93, 8)),
			9756 => std_logic_vector(to_unsigned(24, 8)),
			9757 => std_logic_vector(to_unsigned(122, 8)),
			9758 => std_logic_vector(to_unsigned(207, 8)),
			9759 => std_logic_vector(to_unsigned(89, 8)),
			9760 => std_logic_vector(to_unsigned(48, 8)),
			9761 => std_logic_vector(to_unsigned(163, 8)),
			9762 => std_logic_vector(to_unsigned(29, 8)),
			9763 => std_logic_vector(to_unsigned(84, 8)),
			9764 => std_logic_vector(to_unsigned(248, 8)),
			9765 => std_logic_vector(to_unsigned(41, 8)),
			9766 => std_logic_vector(to_unsigned(91, 8)),
			9767 => std_logic_vector(to_unsigned(203, 8)),
			9768 => std_logic_vector(to_unsigned(14, 8)),
			9769 => std_logic_vector(to_unsigned(244, 8)),
			9770 => std_logic_vector(to_unsigned(37, 8)),
			9771 => std_logic_vector(to_unsigned(90, 8)),
			9772 => std_logic_vector(to_unsigned(211, 8)),
			9773 => std_logic_vector(to_unsigned(37, 8)),
			9774 => std_logic_vector(to_unsigned(8, 8)),
			9775 => std_logic_vector(to_unsigned(104, 8)),
			9776 => std_logic_vector(to_unsigned(225, 8)),
			9777 => std_logic_vector(to_unsigned(167, 8)),
			9778 => std_logic_vector(to_unsigned(151, 8)),
			9779 => std_logic_vector(to_unsigned(203, 8)),
			9780 => std_logic_vector(to_unsigned(246, 8)),
			9781 => std_logic_vector(to_unsigned(147, 8)),
			9782 => std_logic_vector(to_unsigned(158, 8)),
			9783 => std_logic_vector(to_unsigned(145, 8)),
			9784 => std_logic_vector(to_unsigned(153, 8)),
			9785 => std_logic_vector(to_unsigned(197, 8)),
			9786 => std_logic_vector(to_unsigned(46, 8)),
			9787 => std_logic_vector(to_unsigned(115, 8)),
			9788 => std_logic_vector(to_unsigned(82, 8)),
			9789 => std_logic_vector(to_unsigned(15, 8)),
			9790 => std_logic_vector(to_unsigned(25, 8)),
			9791 => std_logic_vector(to_unsigned(131, 8)),
			9792 => std_logic_vector(to_unsigned(20, 8)),
			9793 => std_logic_vector(to_unsigned(230, 8)),
			9794 => std_logic_vector(to_unsigned(227, 8)),
			9795 => std_logic_vector(to_unsigned(152, 8)),
			9796 => std_logic_vector(to_unsigned(94, 8)),
			9797 => std_logic_vector(to_unsigned(34, 8)),
			9798 => std_logic_vector(to_unsigned(159, 8)),
			9799 => std_logic_vector(to_unsigned(112, 8)),
			9800 => std_logic_vector(to_unsigned(134, 8)),
			9801 => std_logic_vector(to_unsigned(210, 8)),
			9802 => std_logic_vector(to_unsigned(204, 8)),
			9803 => std_logic_vector(to_unsigned(145, 8)),
			9804 => std_logic_vector(to_unsigned(139, 8)),
			9805 => std_logic_vector(to_unsigned(144, 8)),
			9806 => std_logic_vector(to_unsigned(65, 8)),
			9807 => std_logic_vector(to_unsigned(165, 8)),
			9808 => std_logic_vector(to_unsigned(194, 8)),
			9809 => std_logic_vector(to_unsigned(246, 8)),
			9810 => std_logic_vector(to_unsigned(186, 8)),
			9811 => std_logic_vector(to_unsigned(94, 8)),
			9812 => std_logic_vector(to_unsigned(61, 8)),
			9813 => std_logic_vector(to_unsigned(142, 8)),
			9814 => std_logic_vector(to_unsigned(240, 8)),
			9815 => std_logic_vector(to_unsigned(3, 8)),
			9816 => std_logic_vector(to_unsigned(170, 8)),
			9817 => std_logic_vector(to_unsigned(184, 8)),
			9818 => std_logic_vector(to_unsigned(83, 8)),
			9819 => std_logic_vector(to_unsigned(222, 8)),
			9820 => std_logic_vector(to_unsigned(73, 8)),
			9821 => std_logic_vector(to_unsigned(77, 8)),
			9822 => std_logic_vector(to_unsigned(70, 8)),
			9823 => std_logic_vector(to_unsigned(253, 8)),
			9824 => std_logic_vector(to_unsigned(189, 8)),
			9825 => std_logic_vector(to_unsigned(111, 8)),
			9826 => std_logic_vector(to_unsigned(190, 8)),
			9827 => std_logic_vector(to_unsigned(233, 8)),
			9828 => std_logic_vector(to_unsigned(170, 8)),
			9829 => std_logic_vector(to_unsigned(213, 8)),
			9830 => std_logic_vector(to_unsigned(103, 8)),
			9831 => std_logic_vector(to_unsigned(68, 8)),
			9832 => std_logic_vector(to_unsigned(97, 8)),
			9833 => std_logic_vector(to_unsigned(31, 8)),
			9834 => std_logic_vector(to_unsigned(214, 8)),
			9835 => std_logic_vector(to_unsigned(129, 8)),
			9836 => std_logic_vector(to_unsigned(219, 8)),
			9837 => std_logic_vector(to_unsigned(161, 8)),
			9838 => std_logic_vector(to_unsigned(38, 8)),
			9839 => std_logic_vector(to_unsigned(105, 8)),
			9840 => std_logic_vector(to_unsigned(37, 8)),
			9841 => std_logic_vector(to_unsigned(119, 8)),
			9842 => std_logic_vector(to_unsigned(231, 8)),
			9843 => std_logic_vector(to_unsigned(193, 8)),
			9844 => std_logic_vector(to_unsigned(226, 8)),
			9845 => std_logic_vector(to_unsigned(212, 8)),
			9846 => std_logic_vector(to_unsigned(17, 8)),
			9847 => std_logic_vector(to_unsigned(171, 8)),
			9848 => std_logic_vector(to_unsigned(122, 8)),
			9849 => std_logic_vector(to_unsigned(121, 8)),
			9850 => std_logic_vector(to_unsigned(91, 8)),
			9851 => std_logic_vector(to_unsigned(224, 8)),
			9852 => std_logic_vector(to_unsigned(233, 8)),
			9853 => std_logic_vector(to_unsigned(8, 8)),
			9854 => std_logic_vector(to_unsigned(211, 8)),
			9855 => std_logic_vector(to_unsigned(151, 8)),
			9856 => std_logic_vector(to_unsigned(252, 8)),
			9857 => std_logic_vector(to_unsigned(23, 8)),
			9858 => std_logic_vector(to_unsigned(149, 8)),
			9859 => std_logic_vector(to_unsigned(226, 8)),
			9860 => std_logic_vector(to_unsigned(119, 8)),
			9861 => std_logic_vector(to_unsigned(37, 8)),
			9862 => std_logic_vector(to_unsigned(139, 8)),
			9863 => std_logic_vector(to_unsigned(213, 8)),
			9864 => std_logic_vector(to_unsigned(171, 8)),
			9865 => std_logic_vector(to_unsigned(222, 8)),
			9866 => std_logic_vector(to_unsigned(42, 8)),
			9867 => std_logic_vector(to_unsigned(37, 8)),
			9868 => std_logic_vector(to_unsigned(182, 8)),
			9869 => std_logic_vector(to_unsigned(175, 8)),
			9870 => std_logic_vector(to_unsigned(149, 8)),
			9871 => std_logic_vector(to_unsigned(12, 8)),
			9872 => std_logic_vector(to_unsigned(62, 8)),
			9873 => std_logic_vector(to_unsigned(78, 8)),
			9874 => std_logic_vector(to_unsigned(72, 8)),
			9875 => std_logic_vector(to_unsigned(147, 8)),
			9876 => std_logic_vector(to_unsigned(200, 8)),
			9877 => std_logic_vector(to_unsigned(171, 8)),
			9878 => std_logic_vector(to_unsigned(197, 8)),
			9879 => std_logic_vector(to_unsigned(236, 8)),
			9880 => std_logic_vector(to_unsigned(69, 8)),
			9881 => std_logic_vector(to_unsigned(250, 8)),
			9882 => std_logic_vector(to_unsigned(182, 8)),
			9883 => std_logic_vector(to_unsigned(51, 8)),
			9884 => std_logic_vector(to_unsigned(150, 8)),
			9885 => std_logic_vector(to_unsigned(7, 8)),
			9886 => std_logic_vector(to_unsigned(184, 8)),
			9887 => std_logic_vector(to_unsigned(8, 8)),
			9888 => std_logic_vector(to_unsigned(202, 8)),
			9889 => std_logic_vector(to_unsigned(9, 8)),
			9890 => std_logic_vector(to_unsigned(35, 8)),
			9891 => std_logic_vector(to_unsigned(185, 8)),
			9892 => std_logic_vector(to_unsigned(155, 8)),
			9893 => std_logic_vector(to_unsigned(158, 8)),
			9894 => std_logic_vector(to_unsigned(37, 8)),
			9895 => std_logic_vector(to_unsigned(209, 8)),
			9896 => std_logic_vector(to_unsigned(35, 8)),
			9897 => std_logic_vector(to_unsigned(42, 8)),
			9898 => std_logic_vector(to_unsigned(108, 8)),
			9899 => std_logic_vector(to_unsigned(127, 8)),
			9900 => std_logic_vector(to_unsigned(140, 8)),
			9901 => std_logic_vector(to_unsigned(71, 8)),
			9902 => std_logic_vector(to_unsigned(206, 8)),
			9903 => std_logic_vector(to_unsigned(219, 8)),
			9904 => std_logic_vector(to_unsigned(228, 8)),
			9905 => std_logic_vector(to_unsigned(25, 8)),
			9906 => std_logic_vector(to_unsigned(203, 8)),
			9907 => std_logic_vector(to_unsigned(51, 8)),
			9908 => std_logic_vector(to_unsigned(173, 8)),
			9909 => std_logic_vector(to_unsigned(253, 8)),
			9910 => std_logic_vector(to_unsigned(11, 8)),
			9911 => std_logic_vector(to_unsigned(157, 8)),
			9912 => std_logic_vector(to_unsigned(216, 8)),
			9913 => std_logic_vector(to_unsigned(235, 8)),
			9914 => std_logic_vector(to_unsigned(53, 8)),
			9915 => std_logic_vector(to_unsigned(193, 8)),
			9916 => std_logic_vector(to_unsigned(25, 8)),
			9917 => std_logic_vector(to_unsigned(207, 8)),
			9918 => std_logic_vector(to_unsigned(249, 8)),
			9919 => std_logic_vector(to_unsigned(56, 8)),
			9920 => std_logic_vector(to_unsigned(3, 8)),
			9921 => std_logic_vector(to_unsigned(12, 8)),
			9922 => std_logic_vector(to_unsigned(240, 8)),
			9923 => std_logic_vector(to_unsigned(215, 8)),
			9924 => std_logic_vector(to_unsigned(50, 8)),
			9925 => std_logic_vector(to_unsigned(209, 8)),
			9926 => std_logic_vector(to_unsigned(61, 8)),
			9927 => std_logic_vector(to_unsigned(104, 8)),
			9928 => std_logic_vector(to_unsigned(242, 8)),
			9929 => std_logic_vector(to_unsigned(90, 8)),
			9930 => std_logic_vector(to_unsigned(153, 8)),
			9931 => std_logic_vector(to_unsigned(37, 8)),
			9932 => std_logic_vector(to_unsigned(85, 8)),
			9933 => std_logic_vector(to_unsigned(226, 8)),
			9934 => std_logic_vector(to_unsigned(70, 8)),
			9935 => std_logic_vector(to_unsigned(46, 8)),
			9936 => std_logic_vector(to_unsigned(73, 8)),
			9937 => std_logic_vector(to_unsigned(171, 8)),
			9938 => std_logic_vector(to_unsigned(242, 8)),
			9939 => std_logic_vector(to_unsigned(2, 8)),
			9940 => std_logic_vector(to_unsigned(204, 8)),
			9941 => std_logic_vector(to_unsigned(87, 8)),
			9942 => std_logic_vector(to_unsigned(45, 8)),
			9943 => std_logic_vector(to_unsigned(44, 8)),
			9944 => std_logic_vector(to_unsigned(58, 8)),
			9945 => std_logic_vector(to_unsigned(89, 8)),
			9946 => std_logic_vector(to_unsigned(4, 8)),
			9947 => std_logic_vector(to_unsigned(212, 8)),
			9948 => std_logic_vector(to_unsigned(221, 8)),
			9949 => std_logic_vector(to_unsigned(241, 8)),
			9950 => std_logic_vector(to_unsigned(107, 8)),
			9951 => std_logic_vector(to_unsigned(202, 8)),
			9952 => std_logic_vector(to_unsigned(61, 8)),
			9953 => std_logic_vector(to_unsigned(255, 8)),
			9954 => std_logic_vector(to_unsigned(212, 8)),
			9955 => std_logic_vector(to_unsigned(136, 8)),
			9956 => std_logic_vector(to_unsigned(206, 8)),
			9957 => std_logic_vector(to_unsigned(184, 8)),
			9958 => std_logic_vector(to_unsigned(241, 8)),
			9959 => std_logic_vector(to_unsigned(43, 8)),
			9960 => std_logic_vector(to_unsigned(108, 8)),
			9961 => std_logic_vector(to_unsigned(36, 8)),
			9962 => std_logic_vector(to_unsigned(47, 8)),
			9963 => std_logic_vector(to_unsigned(217, 8)),
			9964 => std_logic_vector(to_unsigned(127, 8)),
			9965 => std_logic_vector(to_unsigned(200, 8)),
			9966 => std_logic_vector(to_unsigned(0, 8)),
			9967 => std_logic_vector(to_unsigned(150, 8)),
			9968 => std_logic_vector(to_unsigned(252, 8)),
			9969 => std_logic_vector(to_unsigned(69, 8)),
			9970 => std_logic_vector(to_unsigned(39, 8)),
			9971 => std_logic_vector(to_unsigned(57, 8)),
			9972 => std_logic_vector(to_unsigned(220, 8)),
			9973 => std_logic_vector(to_unsigned(209, 8)),
			9974 => std_logic_vector(to_unsigned(16, 8)),
			9975 => std_logic_vector(to_unsigned(182, 8)),
			9976 => std_logic_vector(to_unsigned(169, 8)),
			9977 => std_logic_vector(to_unsigned(110, 8)),
			9978 => std_logic_vector(to_unsigned(237, 8)),
			9979 => std_logic_vector(to_unsigned(7, 8)),
			9980 => std_logic_vector(to_unsigned(179, 8)),
			9981 => std_logic_vector(to_unsigned(99, 8)),
			9982 => std_logic_vector(to_unsigned(16, 8)),
			9983 => std_logic_vector(to_unsigned(89, 8)),
			9984 => std_logic_vector(to_unsigned(142, 8)),
			9985 => std_logic_vector(to_unsigned(84, 8)),
			9986 => std_logic_vector(to_unsigned(86, 8)),
			9987 => std_logic_vector(to_unsigned(95, 8)),
			9988 => std_logic_vector(to_unsigned(116, 8)),
			9989 => std_logic_vector(to_unsigned(74, 8)),
			9990 => std_logic_vector(to_unsigned(146, 8)),
			9991 => std_logic_vector(to_unsigned(7, 8)),
			9992 => std_logic_vector(to_unsigned(65, 8)),
			9993 => std_logic_vector(to_unsigned(8, 8)),
			9994 => std_logic_vector(to_unsigned(213, 8)),
			9995 => std_logic_vector(to_unsigned(87, 8)),
			9996 => std_logic_vector(to_unsigned(56, 8)),
			9997 => std_logic_vector(to_unsigned(16, 8)),
			9998 => std_logic_vector(to_unsigned(61, 8)),
			9999 => std_logic_vector(to_unsigned(224, 8)),
			10000 => std_logic_vector(to_unsigned(73, 8)),
			10001 => std_logic_vector(to_unsigned(234, 8)),
			10002 => std_logic_vector(to_unsigned(85, 8)),
			10003 => std_logic_vector(to_unsigned(156, 8)),
			10004 => std_logic_vector(to_unsigned(105, 8)),
			10005 => std_logic_vector(to_unsigned(36, 8)),
			10006 => std_logic_vector(to_unsigned(48, 8)),
			10007 => std_logic_vector(to_unsigned(139, 8)),
			10008 => std_logic_vector(to_unsigned(130, 8)),
			10009 => std_logic_vector(to_unsigned(175, 8)),
			10010 => std_logic_vector(to_unsigned(9, 8)),
			10011 => std_logic_vector(to_unsigned(26, 8)),
			10012 => std_logic_vector(to_unsigned(217, 8)),
			10013 => std_logic_vector(to_unsigned(97, 8)),
			10014 => std_logic_vector(to_unsigned(1, 8)),
			10015 => std_logic_vector(to_unsigned(16, 8)),
			10016 => std_logic_vector(to_unsigned(165, 8)),
			10017 => std_logic_vector(to_unsigned(84, 8)),
			10018 => std_logic_vector(to_unsigned(84, 8)),
			10019 => std_logic_vector(to_unsigned(41, 8)),
			10020 => std_logic_vector(to_unsigned(67, 8)),
			10021 => std_logic_vector(to_unsigned(182, 8)),
			10022 => std_logic_vector(to_unsigned(149, 8)),
			10023 => std_logic_vector(to_unsigned(88, 8)),
			10024 => std_logic_vector(to_unsigned(254, 8)),
			10025 => std_logic_vector(to_unsigned(230, 8)),
			10026 => std_logic_vector(to_unsigned(29, 8)),
			10027 => std_logic_vector(to_unsigned(45, 8)),
			10028 => std_logic_vector(to_unsigned(36, 8)),
			10029 => std_logic_vector(to_unsigned(204, 8)),
			10030 => std_logic_vector(to_unsigned(134, 8)),
			10031 => std_logic_vector(to_unsigned(95, 8)),
			10032 => std_logic_vector(to_unsigned(201, 8)),
			10033 => std_logic_vector(to_unsigned(229, 8)),
			10034 => std_logic_vector(to_unsigned(19, 8)),
			10035 => std_logic_vector(to_unsigned(167, 8)),
			10036 => std_logic_vector(to_unsigned(67, 8)),
			10037 => std_logic_vector(to_unsigned(111, 8)),
			10038 => std_logic_vector(to_unsigned(70, 8)),
			10039 => std_logic_vector(to_unsigned(250, 8)),
			10040 => std_logic_vector(to_unsigned(121, 8)),
			10041 => std_logic_vector(to_unsigned(216, 8)),
			10042 => std_logic_vector(to_unsigned(130, 8)),
			10043 => std_logic_vector(to_unsigned(95, 8)),
			10044 => std_logic_vector(to_unsigned(121, 8)),
			10045 => std_logic_vector(to_unsigned(153, 8)),
			10046 => std_logic_vector(to_unsigned(9, 8)),
			10047 => std_logic_vector(to_unsigned(216, 8)),
			10048 => std_logic_vector(to_unsigned(7, 8)),
			10049 => std_logic_vector(to_unsigned(47, 8)),
			10050 => std_logic_vector(to_unsigned(44, 8)),
			10051 => std_logic_vector(to_unsigned(56, 8)),
			10052 => std_logic_vector(to_unsigned(147, 8)),
			10053 => std_logic_vector(to_unsigned(124, 8)),
			10054 => std_logic_vector(to_unsigned(13, 8)),
			10055 => std_logic_vector(to_unsigned(115, 8)),
			10056 => std_logic_vector(to_unsigned(210, 8)),
			10057 => std_logic_vector(to_unsigned(255, 8)),
			10058 => std_logic_vector(to_unsigned(162, 8)),
			10059 => std_logic_vector(to_unsigned(252, 8)),
			10060 => std_logic_vector(to_unsigned(214, 8)),
			10061 => std_logic_vector(to_unsigned(110, 8)),
			10062 => std_logic_vector(to_unsigned(100, 8)),
			10063 => std_logic_vector(to_unsigned(64, 8)),
			10064 => std_logic_vector(to_unsigned(76, 8)),
			10065 => std_logic_vector(to_unsigned(0, 8)),
			10066 => std_logic_vector(to_unsigned(232, 8)),
			10067 => std_logic_vector(to_unsigned(115, 8)),
			10068 => std_logic_vector(to_unsigned(71, 8)),
			10069 => std_logic_vector(to_unsigned(223, 8)),
			10070 => std_logic_vector(to_unsigned(148, 8)),
			10071 => std_logic_vector(to_unsigned(25, 8)),
			10072 => std_logic_vector(to_unsigned(21, 8)),
			10073 => std_logic_vector(to_unsigned(61, 8)),
			10074 => std_logic_vector(to_unsigned(253, 8)),
			10075 => std_logic_vector(to_unsigned(213, 8)),
			10076 => std_logic_vector(to_unsigned(54, 8)),
			10077 => std_logic_vector(to_unsigned(195, 8)),
			10078 => std_logic_vector(to_unsigned(14, 8)),
			10079 => std_logic_vector(to_unsigned(186, 8)),
			10080 => std_logic_vector(to_unsigned(9, 8)),
			10081 => std_logic_vector(to_unsigned(171, 8)),
			10082 => std_logic_vector(to_unsigned(37, 8)),
			10083 => std_logic_vector(to_unsigned(45, 8)),
			10084 => std_logic_vector(to_unsigned(195, 8)),
			10085 => std_logic_vector(to_unsigned(112, 8)),
			10086 => std_logic_vector(to_unsigned(73, 8)),
			10087 => std_logic_vector(to_unsigned(147, 8)),
			10088 => std_logic_vector(to_unsigned(57, 8)),
			10089 => std_logic_vector(to_unsigned(220, 8)),
			10090 => std_logic_vector(to_unsigned(45, 8)),
			10091 => std_logic_vector(to_unsigned(63, 8)),
			10092 => std_logic_vector(to_unsigned(215, 8)),
			10093 => std_logic_vector(to_unsigned(248, 8)),
			10094 => std_logic_vector(to_unsigned(242, 8)),
			10095 => std_logic_vector(to_unsigned(138, 8)),
			10096 => std_logic_vector(to_unsigned(72, 8)),
			10097 => std_logic_vector(to_unsigned(106, 8)),
			10098 => std_logic_vector(to_unsigned(246, 8)),
			10099 => std_logic_vector(to_unsigned(166, 8)),
			10100 => std_logic_vector(to_unsigned(6, 8)),
			10101 => std_logic_vector(to_unsigned(75, 8)),
			10102 => std_logic_vector(to_unsigned(51, 8)),
			10103 => std_logic_vector(to_unsigned(16, 8)),
			10104 => std_logic_vector(to_unsigned(184, 8)),
			10105 => std_logic_vector(to_unsigned(84, 8)),
			10106 => std_logic_vector(to_unsigned(193, 8)),
			10107 => std_logic_vector(to_unsigned(104, 8)),
			10108 => std_logic_vector(to_unsigned(246, 8)),
			10109 => std_logic_vector(to_unsigned(14, 8)),
			10110 => std_logic_vector(to_unsigned(98, 8)),
			10111 => std_logic_vector(to_unsigned(208, 8)),
			10112 => std_logic_vector(to_unsigned(119, 8)),
			10113 => std_logic_vector(to_unsigned(161, 8)),
			10114 => std_logic_vector(to_unsigned(169, 8)),
			10115 => std_logic_vector(to_unsigned(239, 8)),
			10116 => std_logic_vector(to_unsigned(11, 8)),
			10117 => std_logic_vector(to_unsigned(51, 8)),
			10118 => std_logic_vector(to_unsigned(168, 8)),
			10119 => std_logic_vector(to_unsigned(101, 8)),
			10120 => std_logic_vector(to_unsigned(212, 8)),
			10121 => std_logic_vector(to_unsigned(138, 8)),
			10122 => std_logic_vector(to_unsigned(48, 8)),
			10123 => std_logic_vector(to_unsigned(0, 8)),
			10124 => std_logic_vector(to_unsigned(232, 8)),
			10125 => std_logic_vector(to_unsigned(98, 8)),
			10126 => std_logic_vector(to_unsigned(199, 8)),
			10127 => std_logic_vector(to_unsigned(147, 8)),
			10128 => std_logic_vector(to_unsigned(243, 8)),
			10129 => std_logic_vector(to_unsigned(120, 8)),
			10130 => std_logic_vector(to_unsigned(154, 8)),
			10131 => std_logic_vector(to_unsigned(182, 8)),
			10132 => std_logic_vector(to_unsigned(223, 8)),
			10133 => std_logic_vector(to_unsigned(213, 8)),
			10134 => std_logic_vector(to_unsigned(137, 8)),
			10135 => std_logic_vector(to_unsigned(105, 8)),
			10136 => std_logic_vector(to_unsigned(24, 8)),
			10137 => std_logic_vector(to_unsigned(76, 8)),
			10138 => std_logic_vector(to_unsigned(60, 8)),
			10139 => std_logic_vector(to_unsigned(43, 8)),
			10140 => std_logic_vector(to_unsigned(61, 8)),
			10141 => std_logic_vector(to_unsigned(109, 8)),
			10142 => std_logic_vector(to_unsigned(64, 8)),
			10143 => std_logic_vector(to_unsigned(212, 8)),
			10144 => std_logic_vector(to_unsigned(80, 8)),
			10145 => std_logic_vector(to_unsigned(89, 8)),
			10146 => std_logic_vector(to_unsigned(87, 8)),
			10147 => std_logic_vector(to_unsigned(238, 8)),
			10148 => std_logic_vector(to_unsigned(27, 8)),
			10149 => std_logic_vector(to_unsigned(214, 8)),
			10150 => std_logic_vector(to_unsigned(205, 8)),
			10151 => std_logic_vector(to_unsigned(43, 8)),
			10152 => std_logic_vector(to_unsigned(241, 8)),
			10153 => std_logic_vector(to_unsigned(91, 8)),
			10154 => std_logic_vector(to_unsigned(15, 8)),
			10155 => std_logic_vector(to_unsigned(109, 8)),
			10156 => std_logic_vector(to_unsigned(128, 8)),
			10157 => std_logic_vector(to_unsigned(139, 8)),
			10158 => std_logic_vector(to_unsigned(132, 8)),
			10159 => std_logic_vector(to_unsigned(22, 8)),
			10160 => std_logic_vector(to_unsigned(56, 8)),
			10161 => std_logic_vector(to_unsigned(208, 8)),
			10162 => std_logic_vector(to_unsigned(42, 8)),
			10163 => std_logic_vector(to_unsigned(192, 8)),
			10164 => std_logic_vector(to_unsigned(88, 8)),
			10165 => std_logic_vector(to_unsigned(129, 8)),
			10166 => std_logic_vector(to_unsigned(70, 8)),
			10167 => std_logic_vector(to_unsigned(162, 8)),
			10168 => std_logic_vector(to_unsigned(72, 8)),
			10169 => std_logic_vector(to_unsigned(246, 8)),
			10170 => std_logic_vector(to_unsigned(243, 8)),
			10171 => std_logic_vector(to_unsigned(185, 8)),
			10172 => std_logic_vector(to_unsigned(30, 8)),
			10173 => std_logic_vector(to_unsigned(82, 8)),
			10174 => std_logic_vector(to_unsigned(19, 8)),
			10175 => std_logic_vector(to_unsigned(134, 8)),
			10176 => std_logic_vector(to_unsigned(53, 8)),
			10177 => std_logic_vector(to_unsigned(54, 8)),
			10178 => std_logic_vector(to_unsigned(17, 8)),
			10179 => std_logic_vector(to_unsigned(163, 8)),
			10180 => std_logic_vector(to_unsigned(229, 8)),
			10181 => std_logic_vector(to_unsigned(233, 8)),
			10182 => std_logic_vector(to_unsigned(68, 8)),
			10183 => std_logic_vector(to_unsigned(179, 8)),
			10184 => std_logic_vector(to_unsigned(159, 8)),
			10185 => std_logic_vector(to_unsigned(23, 8)),
			10186 => std_logic_vector(to_unsigned(100, 8)),
			10187 => std_logic_vector(to_unsigned(13, 8)),
			10188 => std_logic_vector(to_unsigned(170, 8)),
			10189 => std_logic_vector(to_unsigned(167, 8)),
			10190 => std_logic_vector(to_unsigned(177, 8)),
			10191 => std_logic_vector(to_unsigned(117, 8)),
			10192 => std_logic_vector(to_unsigned(132, 8)),
			10193 => std_logic_vector(to_unsigned(15, 8)),
			10194 => std_logic_vector(to_unsigned(97, 8)),
			10195 => std_logic_vector(to_unsigned(140, 8)),
			10196 => std_logic_vector(to_unsigned(125, 8)),
			10197 => std_logic_vector(to_unsigned(7, 8)),
			10198 => std_logic_vector(to_unsigned(221, 8)),
			10199 => std_logic_vector(to_unsigned(124, 8)),
			10200 => std_logic_vector(to_unsigned(151, 8)),
			10201 => std_logic_vector(to_unsigned(64, 8)),
			10202 => std_logic_vector(to_unsigned(156, 8)),
			10203 => std_logic_vector(to_unsigned(204, 8)),
			10204 => std_logic_vector(to_unsigned(109, 8)),
			10205 => std_logic_vector(to_unsigned(43, 8)),
			10206 => std_logic_vector(to_unsigned(31, 8)),
			10207 => std_logic_vector(to_unsigned(205, 8)),
			10208 => std_logic_vector(to_unsigned(89, 8)),
			10209 => std_logic_vector(to_unsigned(172, 8)),
			10210 => std_logic_vector(to_unsigned(144, 8)),
			10211 => std_logic_vector(to_unsigned(8, 8)),
			10212 => std_logic_vector(to_unsigned(198, 8)),
			10213 => std_logic_vector(to_unsigned(172, 8)),
			10214 => std_logic_vector(to_unsigned(239, 8)),
			10215 => std_logic_vector(to_unsigned(2, 8)),
			10216 => std_logic_vector(to_unsigned(187, 8)),
			10217 => std_logic_vector(to_unsigned(130, 8)),
			10218 => std_logic_vector(to_unsigned(140, 8)),
			10219 => std_logic_vector(to_unsigned(180, 8)),
			10220 => std_logic_vector(to_unsigned(33, 8)),
			10221 => std_logic_vector(to_unsigned(198, 8)),
			10222 => std_logic_vector(to_unsigned(82, 8)),
			10223 => std_logic_vector(to_unsigned(3, 8)),
			10224 => std_logic_vector(to_unsigned(214, 8)),
			10225 => std_logic_vector(to_unsigned(59, 8)),
			10226 => std_logic_vector(to_unsigned(94, 8)),
			10227 => std_logic_vector(to_unsigned(168, 8)),
			10228 => std_logic_vector(to_unsigned(226, 8)),
			10229 => std_logic_vector(to_unsigned(198, 8)),
			10230 => std_logic_vector(to_unsigned(94, 8)),
			10231 => std_logic_vector(to_unsigned(100, 8)),
			10232 => std_logic_vector(to_unsigned(122, 8)),
			10233 => std_logic_vector(to_unsigned(94, 8)),
			10234 => std_logic_vector(to_unsigned(31, 8)),
			10235 => std_logic_vector(to_unsigned(175, 8)),
			10236 => std_logic_vector(to_unsigned(48, 8)),
			10237 => std_logic_vector(to_unsigned(18, 8)),
			10238 => std_logic_vector(to_unsigned(236, 8)),
			10239 => std_logic_vector(to_unsigned(209, 8)),
			10240 => std_logic_vector(to_unsigned(61, 8)),
			10241 => std_logic_vector(to_unsigned(38, 8)),
			10242 => std_logic_vector(to_unsigned(148, 8)),
			10243 => std_logic_vector(to_unsigned(252, 8)),
			10244 => std_logic_vector(to_unsigned(44, 8)),
			10245 => std_logic_vector(to_unsigned(249, 8)),
			10246 => std_logic_vector(to_unsigned(99, 8)),
			10247 => std_logic_vector(to_unsigned(249, 8)),
			10248 => std_logic_vector(to_unsigned(212, 8)),
			10249 => std_logic_vector(to_unsigned(88, 8)),
			10250 => std_logic_vector(to_unsigned(254, 8)),
			10251 => std_logic_vector(to_unsigned(49, 8)),
			10252 => std_logic_vector(to_unsigned(174, 8)),
			10253 => std_logic_vector(to_unsigned(230, 8)),
			10254 => std_logic_vector(to_unsigned(39, 8)),
			10255 => std_logic_vector(to_unsigned(25, 8)),
			10256 => std_logic_vector(to_unsigned(143, 8)),
			10257 => std_logic_vector(to_unsigned(4, 8)),
			10258 => std_logic_vector(to_unsigned(219, 8)),
			10259 => std_logic_vector(to_unsigned(180, 8)),
			10260 => std_logic_vector(to_unsigned(228, 8)),
			10261 => std_logic_vector(to_unsigned(85, 8)),
			10262 => std_logic_vector(to_unsigned(5, 8)),
			10263 => std_logic_vector(to_unsigned(167, 8)),
			10264 => std_logic_vector(to_unsigned(240, 8)),
			10265 => std_logic_vector(to_unsigned(204, 8)),
			10266 => std_logic_vector(to_unsigned(172, 8)),
			10267 => std_logic_vector(to_unsigned(251, 8)),
			10268 => std_logic_vector(to_unsigned(86, 8)),
			10269 => std_logic_vector(to_unsigned(197, 8)),
			10270 => std_logic_vector(to_unsigned(80, 8)),
			10271 => std_logic_vector(to_unsigned(247, 8)),
			10272 => std_logic_vector(to_unsigned(216, 8)),
			10273 => std_logic_vector(to_unsigned(154, 8)),
			10274 => std_logic_vector(to_unsigned(96, 8)),
			10275 => std_logic_vector(to_unsigned(217, 8)),
			10276 => std_logic_vector(to_unsigned(77, 8)),
			10277 => std_logic_vector(to_unsigned(19, 8)),
			10278 => std_logic_vector(to_unsigned(180, 8)),
			10279 => std_logic_vector(to_unsigned(102, 8)),
			10280 => std_logic_vector(to_unsigned(201, 8)),
			10281 => std_logic_vector(to_unsigned(141, 8)),
			10282 => std_logic_vector(to_unsigned(225, 8)),
			10283 => std_logic_vector(to_unsigned(115, 8)),
			10284 => std_logic_vector(to_unsigned(34, 8)),
			10285 => std_logic_vector(to_unsigned(87, 8)),
			10286 => std_logic_vector(to_unsigned(220, 8)),
			10287 => std_logic_vector(to_unsigned(223, 8)),
			10288 => std_logic_vector(to_unsigned(96, 8)),
			10289 => std_logic_vector(to_unsigned(0, 8)),
			10290 => std_logic_vector(to_unsigned(204, 8)),
			10291 => std_logic_vector(to_unsigned(63, 8)),
			10292 => std_logic_vector(to_unsigned(116, 8)),
			10293 => std_logic_vector(to_unsigned(67, 8)),
			10294 => std_logic_vector(to_unsigned(158, 8)),
			10295 => std_logic_vector(to_unsigned(71, 8)),
			10296 => std_logic_vector(to_unsigned(49, 8)),
			10297 => std_logic_vector(to_unsigned(159, 8)),
			10298 => std_logic_vector(to_unsigned(105, 8)),
			10299 => std_logic_vector(to_unsigned(23, 8)),
			10300 => std_logic_vector(to_unsigned(189, 8)),
			10301 => std_logic_vector(to_unsigned(207, 8)),
			10302 => std_logic_vector(to_unsigned(108, 8)),
			10303 => std_logic_vector(to_unsigned(95, 8)),
			10304 => std_logic_vector(to_unsigned(124, 8)),
			10305 => std_logic_vector(to_unsigned(72, 8)),
			10306 => std_logic_vector(to_unsigned(18, 8)),
			10307 => std_logic_vector(to_unsigned(119, 8)),
			10308 => std_logic_vector(to_unsigned(104, 8)),
			10309 => std_logic_vector(to_unsigned(91, 8)),
			10310 => std_logic_vector(to_unsigned(206, 8)),
			10311 => std_logic_vector(to_unsigned(70, 8)),
			10312 => std_logic_vector(to_unsigned(91, 8)),
			10313 => std_logic_vector(to_unsigned(66, 8)),
			10314 => std_logic_vector(to_unsigned(69, 8)),
			10315 => std_logic_vector(to_unsigned(160, 8)),
			10316 => std_logic_vector(to_unsigned(100, 8)),
			10317 => std_logic_vector(to_unsigned(7, 8)),
			10318 => std_logic_vector(to_unsigned(17, 8)),
			10319 => std_logic_vector(to_unsigned(140, 8)),
			10320 => std_logic_vector(to_unsigned(185, 8)),
			10321 => std_logic_vector(to_unsigned(49, 8)),
			10322 => std_logic_vector(to_unsigned(87, 8)),
			10323 => std_logic_vector(to_unsigned(111, 8)),
			10324 => std_logic_vector(to_unsigned(151, 8)),
			10325 => std_logic_vector(to_unsigned(123, 8)),
			10326 => std_logic_vector(to_unsigned(33, 8)),
			10327 => std_logic_vector(to_unsigned(165, 8)),
			10328 => std_logic_vector(to_unsigned(170, 8)),
			10329 => std_logic_vector(to_unsigned(220, 8)),
			10330 => std_logic_vector(to_unsigned(14, 8)),
			10331 => std_logic_vector(to_unsigned(33, 8)),
			10332 => std_logic_vector(to_unsigned(25, 8)),
			10333 => std_logic_vector(to_unsigned(38, 8)),
			10334 => std_logic_vector(to_unsigned(124, 8)),
			10335 => std_logic_vector(to_unsigned(109, 8)),
			10336 => std_logic_vector(to_unsigned(129, 8)),
			10337 => std_logic_vector(to_unsigned(153, 8)),
			10338 => std_logic_vector(to_unsigned(101, 8)),
			10339 => std_logic_vector(to_unsigned(69, 8)),
			10340 => std_logic_vector(to_unsigned(191, 8)),
			10341 => std_logic_vector(to_unsigned(161, 8)),
			10342 => std_logic_vector(to_unsigned(123, 8)),
			10343 => std_logic_vector(to_unsigned(166, 8)),
			10344 => std_logic_vector(to_unsigned(92, 8)),
			10345 => std_logic_vector(to_unsigned(188, 8)),
			10346 => std_logic_vector(to_unsigned(39, 8)),
			10347 => std_logic_vector(to_unsigned(210, 8)),
			10348 => std_logic_vector(to_unsigned(136, 8)),
			10349 => std_logic_vector(to_unsigned(108, 8)),
			10350 => std_logic_vector(to_unsigned(118, 8)),
			10351 => std_logic_vector(to_unsigned(109, 8)),
			10352 => std_logic_vector(to_unsigned(26, 8)),
			10353 => std_logic_vector(to_unsigned(157, 8)),
			10354 => std_logic_vector(to_unsigned(25, 8)),
			10355 => std_logic_vector(to_unsigned(169, 8)),
			10356 => std_logic_vector(to_unsigned(50, 8)),
			10357 => std_logic_vector(to_unsigned(123, 8)),
			10358 => std_logic_vector(to_unsigned(145, 8)),
			10359 => std_logic_vector(to_unsigned(219, 8)),
			10360 => std_logic_vector(to_unsigned(67, 8)),
			10361 => std_logic_vector(to_unsigned(123, 8)),
			10362 => std_logic_vector(to_unsigned(34, 8)),
			10363 => std_logic_vector(to_unsigned(186, 8)),
			10364 => std_logic_vector(to_unsigned(122, 8)),
			10365 => std_logic_vector(to_unsigned(97, 8)),
			10366 => std_logic_vector(to_unsigned(57, 8)),
			10367 => std_logic_vector(to_unsigned(39, 8)),
			10368 => std_logic_vector(to_unsigned(21, 8)),
			10369 => std_logic_vector(to_unsigned(118, 8)),
			10370 => std_logic_vector(to_unsigned(157, 8)),
			10371 => std_logic_vector(to_unsigned(49, 8)),
			10372 => std_logic_vector(to_unsigned(78, 8)),
			10373 => std_logic_vector(to_unsigned(140, 8)),
			10374 => std_logic_vector(to_unsigned(19, 8)),
			10375 => std_logic_vector(to_unsigned(179, 8)),
			10376 => std_logic_vector(to_unsigned(247, 8)),
			10377 => std_logic_vector(to_unsigned(42, 8)),
			10378 => std_logic_vector(to_unsigned(79, 8)),
			10379 => std_logic_vector(to_unsigned(153, 8)),
			10380 => std_logic_vector(to_unsigned(199, 8)),
			10381 => std_logic_vector(to_unsigned(31, 8)),
			10382 => std_logic_vector(to_unsigned(137, 8)),
			10383 => std_logic_vector(to_unsigned(146, 8)),
			10384 => std_logic_vector(to_unsigned(96, 8)),
			10385 => std_logic_vector(to_unsigned(140, 8)),
			10386 => std_logic_vector(to_unsigned(58, 8)),
			10387 => std_logic_vector(to_unsigned(119, 8)),
			10388 => std_logic_vector(to_unsigned(66, 8)),
			10389 => std_logic_vector(to_unsigned(229, 8)),
			10390 => std_logic_vector(to_unsigned(142, 8)),
			10391 => std_logic_vector(to_unsigned(19, 8)),
			10392 => std_logic_vector(to_unsigned(158, 8)),
			10393 => std_logic_vector(to_unsigned(10, 8)),
			10394 => std_logic_vector(to_unsigned(247, 8)),
			10395 => std_logic_vector(to_unsigned(84, 8)),
			10396 => std_logic_vector(to_unsigned(140, 8)),
			10397 => std_logic_vector(to_unsigned(85, 8)),
			10398 => std_logic_vector(to_unsigned(199, 8)),
			10399 => std_logic_vector(to_unsigned(151, 8)),
			10400 => std_logic_vector(to_unsigned(232, 8)),
			10401 => std_logic_vector(to_unsigned(22, 8)),
			10402 => std_logic_vector(to_unsigned(192, 8)),
			10403 => std_logic_vector(to_unsigned(184, 8)),
			10404 => std_logic_vector(to_unsigned(233, 8)),
			10405 => std_logic_vector(to_unsigned(13, 8)),
			10406 => std_logic_vector(to_unsigned(44, 8)),
			10407 => std_logic_vector(to_unsigned(82, 8)),
			10408 => std_logic_vector(to_unsigned(249, 8)),
			10409 => std_logic_vector(to_unsigned(111, 8)),
			10410 => std_logic_vector(to_unsigned(245, 8)),
			10411 => std_logic_vector(to_unsigned(121, 8)),
			10412 => std_logic_vector(to_unsigned(49, 8)),
			10413 => std_logic_vector(to_unsigned(167, 8)),
			10414 => std_logic_vector(to_unsigned(254, 8)),
			10415 => std_logic_vector(to_unsigned(220, 8)),
			10416 => std_logic_vector(to_unsigned(154, 8)),
			10417 => std_logic_vector(to_unsigned(27, 8)),
			10418 => std_logic_vector(to_unsigned(204, 8)),
			10419 => std_logic_vector(to_unsigned(190, 8)),
			10420 => std_logic_vector(to_unsigned(65, 8)),
			10421 => std_logic_vector(to_unsigned(38, 8)),
			10422 => std_logic_vector(to_unsigned(6, 8)),
			10423 => std_logic_vector(to_unsigned(67, 8)),
			10424 => std_logic_vector(to_unsigned(58, 8)),
			10425 => std_logic_vector(to_unsigned(108, 8)),
			10426 => std_logic_vector(to_unsigned(229, 8)),
			10427 => std_logic_vector(to_unsigned(120, 8)),
			10428 => std_logic_vector(to_unsigned(229, 8)),
			10429 => std_logic_vector(to_unsigned(154, 8)),
			10430 => std_logic_vector(to_unsigned(65, 8)),
			10431 => std_logic_vector(to_unsigned(23, 8)),
			10432 => std_logic_vector(to_unsigned(51, 8)),
			10433 => std_logic_vector(to_unsigned(104, 8)),
			10434 => std_logic_vector(to_unsigned(254, 8)),
			10435 => std_logic_vector(to_unsigned(77, 8)),
			10436 => std_logic_vector(to_unsigned(89, 8)),
			10437 => std_logic_vector(to_unsigned(240, 8)),
			10438 => std_logic_vector(to_unsigned(38, 8)),
			10439 => std_logic_vector(to_unsigned(184, 8)),
			10440 => std_logic_vector(to_unsigned(196, 8)),
			10441 => std_logic_vector(to_unsigned(174, 8)),
			10442 => std_logic_vector(to_unsigned(54, 8)),
			10443 => std_logic_vector(to_unsigned(128, 8)),
			10444 => std_logic_vector(to_unsigned(0, 8)),
			10445 => std_logic_vector(to_unsigned(9, 8)),
			10446 => std_logic_vector(to_unsigned(121, 8)),
			10447 => std_logic_vector(to_unsigned(123, 8)),
			10448 => std_logic_vector(to_unsigned(88, 8)),
			10449 => std_logic_vector(to_unsigned(162, 8)),
			10450 => std_logic_vector(to_unsigned(45, 8)),
			10451 => std_logic_vector(to_unsigned(3, 8)),
			10452 => std_logic_vector(to_unsigned(251, 8)),
			10453 => std_logic_vector(to_unsigned(185, 8)),
			10454 => std_logic_vector(to_unsigned(67, 8)),
			10455 => std_logic_vector(to_unsigned(178, 8)),
			10456 => std_logic_vector(to_unsigned(224, 8)),
			10457 => std_logic_vector(to_unsigned(185, 8)),
			10458 => std_logic_vector(to_unsigned(136, 8)),
			10459 => std_logic_vector(to_unsigned(240, 8)),
			10460 => std_logic_vector(to_unsigned(250, 8)),
			10461 => std_logic_vector(to_unsigned(107, 8)),
			10462 => std_logic_vector(to_unsigned(214, 8)),
			10463 => std_logic_vector(to_unsigned(45, 8)),
			10464 => std_logic_vector(to_unsigned(9, 8)),
			10465 => std_logic_vector(to_unsigned(148, 8)),
			10466 => std_logic_vector(to_unsigned(142, 8)),
			10467 => std_logic_vector(to_unsigned(249, 8)),
			10468 => std_logic_vector(to_unsigned(218, 8)),
			10469 => std_logic_vector(to_unsigned(152, 8)),
			10470 => std_logic_vector(to_unsigned(94, 8)),
			10471 => std_logic_vector(to_unsigned(8, 8)),
			10472 => std_logic_vector(to_unsigned(170, 8)),
			10473 => std_logic_vector(to_unsigned(54, 8)),
			10474 => std_logic_vector(to_unsigned(190, 8)),
			10475 => std_logic_vector(to_unsigned(239, 8)),
			10476 => std_logic_vector(to_unsigned(211, 8)),
			10477 => std_logic_vector(to_unsigned(57, 8)),
			10478 => std_logic_vector(to_unsigned(45, 8)),
			10479 => std_logic_vector(to_unsigned(252, 8)),
			10480 => std_logic_vector(to_unsigned(182, 8)),
			10481 => std_logic_vector(to_unsigned(54, 8)),
			10482 => std_logic_vector(to_unsigned(45, 8)),
			10483 => std_logic_vector(to_unsigned(72, 8)),
			10484 => std_logic_vector(to_unsigned(61, 8)),
			10485 => std_logic_vector(to_unsigned(217, 8)),
			10486 => std_logic_vector(to_unsigned(10, 8)),
			10487 => std_logic_vector(to_unsigned(144, 8)),
			10488 => std_logic_vector(to_unsigned(106, 8)),
			10489 => std_logic_vector(to_unsigned(195, 8)),
			10490 => std_logic_vector(to_unsigned(11, 8)),
			10491 => std_logic_vector(to_unsigned(217, 8)),
			10492 => std_logic_vector(to_unsigned(228, 8)),
			10493 => std_logic_vector(to_unsigned(246, 8)),
			10494 => std_logic_vector(to_unsigned(126, 8)),
			10495 => std_logic_vector(to_unsigned(39, 8)),
			10496 => std_logic_vector(to_unsigned(214, 8)),
			10497 => std_logic_vector(to_unsigned(82, 8)),
			10498 => std_logic_vector(to_unsigned(31, 8)),
			10499 => std_logic_vector(to_unsigned(227, 8)),
			10500 => std_logic_vector(to_unsigned(61, 8)),
			10501 => std_logic_vector(to_unsigned(165, 8)),
			10502 => std_logic_vector(to_unsigned(208, 8)),
			10503 => std_logic_vector(to_unsigned(104, 8)),
			10504 => std_logic_vector(to_unsigned(117, 8)),
			10505 => std_logic_vector(to_unsigned(96, 8)),
			10506 => std_logic_vector(to_unsigned(118, 8)),
			10507 => std_logic_vector(to_unsigned(36, 8)),
			10508 => std_logic_vector(to_unsigned(72, 8)),
			10509 => std_logic_vector(to_unsigned(119, 8)),
			10510 => std_logic_vector(to_unsigned(251, 8)),
			10511 => std_logic_vector(to_unsigned(76, 8)),
			10512 => std_logic_vector(to_unsigned(24, 8)),
			10513 => std_logic_vector(to_unsigned(26, 8)),
			10514 => std_logic_vector(to_unsigned(47, 8)),
			10515 => std_logic_vector(to_unsigned(233, 8)),
			10516 => std_logic_vector(to_unsigned(155, 8)),
			10517 => std_logic_vector(to_unsigned(195, 8)),
			10518 => std_logic_vector(to_unsigned(114, 8)),
			10519 => std_logic_vector(to_unsigned(226, 8)),
			10520 => std_logic_vector(to_unsigned(250, 8)),
			10521 => std_logic_vector(to_unsigned(107, 8)),
			10522 => std_logic_vector(to_unsigned(58, 8)),
			10523 => std_logic_vector(to_unsigned(59, 8)),
			10524 => std_logic_vector(to_unsigned(184, 8)),
			10525 => std_logic_vector(to_unsigned(67, 8)),
			10526 => std_logic_vector(to_unsigned(97, 8)),
			10527 => std_logic_vector(to_unsigned(135, 8)),
			10528 => std_logic_vector(to_unsigned(10, 8)),
			10529 => std_logic_vector(to_unsigned(98, 8)),
			10530 => std_logic_vector(to_unsigned(33, 8)),
			10531 => std_logic_vector(to_unsigned(71, 8)),
			10532 => std_logic_vector(to_unsigned(30, 8)),
			10533 => std_logic_vector(to_unsigned(211, 8)),
			10534 => std_logic_vector(to_unsigned(230, 8)),
			10535 => std_logic_vector(to_unsigned(82, 8)),
			10536 => std_logic_vector(to_unsigned(54, 8)),
			10537 => std_logic_vector(to_unsigned(49, 8)),
			10538 => std_logic_vector(to_unsigned(22, 8)),
			10539 => std_logic_vector(to_unsigned(199, 8)),
			10540 => std_logic_vector(to_unsigned(220, 8)),
			10541 => std_logic_vector(to_unsigned(192, 8)),
			10542 => std_logic_vector(to_unsigned(222, 8)),
			10543 => std_logic_vector(to_unsigned(163, 8)),
			10544 => std_logic_vector(to_unsigned(69, 8)),
			10545 => std_logic_vector(to_unsigned(31, 8)),
			10546 => std_logic_vector(to_unsigned(150, 8)),
			10547 => std_logic_vector(to_unsigned(25, 8)),
			10548 => std_logic_vector(to_unsigned(39, 8)),
			10549 => std_logic_vector(to_unsigned(195, 8)),
			10550 => std_logic_vector(to_unsigned(96, 8)),
			10551 => std_logic_vector(to_unsigned(230, 8)),
			10552 => std_logic_vector(to_unsigned(20, 8)),
			10553 => std_logic_vector(to_unsigned(1, 8)),
			10554 => std_logic_vector(to_unsigned(221, 8)),
			10555 => std_logic_vector(to_unsigned(238, 8)),
			10556 => std_logic_vector(to_unsigned(86, 8)),
			10557 => std_logic_vector(to_unsigned(112, 8)),
			10558 => std_logic_vector(to_unsigned(179, 8)),
			10559 => std_logic_vector(to_unsigned(190, 8)),
			10560 => std_logic_vector(to_unsigned(105, 8)),
			10561 => std_logic_vector(to_unsigned(149, 8)),
			10562 => std_logic_vector(to_unsigned(191, 8)),
			10563 => std_logic_vector(to_unsigned(93, 8)),
			10564 => std_logic_vector(to_unsigned(55, 8)),
			10565 => std_logic_vector(to_unsigned(27, 8)),
			10566 => std_logic_vector(to_unsigned(49, 8)),
			10567 => std_logic_vector(to_unsigned(184, 8)),
			10568 => std_logic_vector(to_unsigned(177, 8)),
			10569 => std_logic_vector(to_unsigned(143, 8)),
			10570 => std_logic_vector(to_unsigned(240, 8)),
			10571 => std_logic_vector(to_unsigned(40, 8)),
			10572 => std_logic_vector(to_unsigned(3, 8)),
			10573 => std_logic_vector(to_unsigned(139, 8)),
			10574 => std_logic_vector(to_unsigned(18, 8)),
			10575 => std_logic_vector(to_unsigned(38, 8)),
			10576 => std_logic_vector(to_unsigned(181, 8)),
			10577 => std_logic_vector(to_unsigned(165, 8)),
			10578 => std_logic_vector(to_unsigned(74, 8)),
			10579 => std_logic_vector(to_unsigned(205, 8)),
			10580 => std_logic_vector(to_unsigned(13, 8)),
			10581 => std_logic_vector(to_unsigned(77, 8)),
			10582 => std_logic_vector(to_unsigned(46, 8)),
			10583 => std_logic_vector(to_unsigned(38, 8)),
			10584 => std_logic_vector(to_unsigned(86, 8)),
			10585 => std_logic_vector(to_unsigned(188, 8)),
			10586 => std_logic_vector(to_unsigned(73, 8)),
			10587 => std_logic_vector(to_unsigned(182, 8)),
			10588 => std_logic_vector(to_unsigned(223, 8)),
			10589 => std_logic_vector(to_unsigned(190, 8)),
			10590 => std_logic_vector(to_unsigned(87, 8)),
			10591 => std_logic_vector(to_unsigned(18, 8)),
			10592 => std_logic_vector(to_unsigned(61, 8)),
			10593 => std_logic_vector(to_unsigned(102, 8)),
			10594 => std_logic_vector(to_unsigned(72, 8)),
			10595 => std_logic_vector(to_unsigned(210, 8)),
			10596 => std_logic_vector(to_unsigned(167, 8)),
			10597 => std_logic_vector(to_unsigned(65, 8)),
			10598 => std_logic_vector(to_unsigned(2, 8)),
			10599 => std_logic_vector(to_unsigned(98, 8)),
			10600 => std_logic_vector(to_unsigned(13, 8)),
			10601 => std_logic_vector(to_unsigned(22, 8)),
			10602 => std_logic_vector(to_unsigned(147, 8)),
			10603 => std_logic_vector(to_unsigned(87, 8)),
			10604 => std_logic_vector(to_unsigned(81, 8)),
			10605 => std_logic_vector(to_unsigned(157, 8)),
			10606 => std_logic_vector(to_unsigned(175, 8)),
			10607 => std_logic_vector(to_unsigned(99, 8)),
			10608 => std_logic_vector(to_unsigned(230, 8)),
			10609 => std_logic_vector(to_unsigned(222, 8)),
			10610 => std_logic_vector(to_unsigned(97, 8)),
			10611 => std_logic_vector(to_unsigned(5, 8)),
			10612 => std_logic_vector(to_unsigned(130, 8)),
			10613 => std_logic_vector(to_unsigned(212, 8)),
			10614 => std_logic_vector(to_unsigned(217, 8)),
			10615 => std_logic_vector(to_unsigned(186, 8)),
			10616 => std_logic_vector(to_unsigned(0, 8)),
			10617 => std_logic_vector(to_unsigned(14, 8)),
			10618 => std_logic_vector(to_unsigned(155, 8)),
			10619 => std_logic_vector(to_unsigned(255, 8)),
			10620 => std_logic_vector(to_unsigned(158, 8)),
			10621 => std_logic_vector(to_unsigned(108, 8)),
			10622 => std_logic_vector(to_unsigned(53, 8)),
			10623 => std_logic_vector(to_unsigned(200, 8)),
			10624 => std_logic_vector(to_unsigned(92, 8)),
			10625 => std_logic_vector(to_unsigned(166, 8)),
			10626 => std_logic_vector(to_unsigned(121, 8)),
			10627 => std_logic_vector(to_unsigned(246, 8)),
			10628 => std_logic_vector(to_unsigned(137, 8)),
			10629 => std_logic_vector(to_unsigned(147, 8)),
			10630 => std_logic_vector(to_unsigned(21, 8)),
			10631 => std_logic_vector(to_unsigned(102, 8)),
			10632 => std_logic_vector(to_unsigned(134, 8)),
			10633 => std_logic_vector(to_unsigned(9, 8)),
			10634 => std_logic_vector(to_unsigned(125, 8)),
			10635 => std_logic_vector(to_unsigned(198, 8)),
			10636 => std_logic_vector(to_unsigned(247, 8)),
			10637 => std_logic_vector(to_unsigned(10, 8)),
			10638 => std_logic_vector(to_unsigned(78, 8)),
			10639 => std_logic_vector(to_unsigned(108, 8)),
			10640 => std_logic_vector(to_unsigned(161, 8)),
			10641 => std_logic_vector(to_unsigned(69, 8)),
			10642 => std_logic_vector(to_unsigned(0, 8)),
			10643 => std_logic_vector(to_unsigned(248, 8)),
			10644 => std_logic_vector(to_unsigned(60, 8)),
			10645 => std_logic_vector(to_unsigned(30, 8)),
			10646 => std_logic_vector(to_unsigned(181, 8)),
			10647 => std_logic_vector(to_unsigned(119, 8)),
			10648 => std_logic_vector(to_unsigned(147, 8)),
			10649 => std_logic_vector(to_unsigned(159, 8)),
			10650 => std_logic_vector(to_unsigned(66, 8)),
			10651 => std_logic_vector(to_unsigned(17, 8)),
			10652 => std_logic_vector(to_unsigned(129, 8)),
			10653 => std_logic_vector(to_unsigned(184, 8)),
			10654 => std_logic_vector(to_unsigned(72, 8)),
			10655 => std_logic_vector(to_unsigned(211, 8)),
			10656 => std_logic_vector(to_unsigned(171, 8)),
			10657 => std_logic_vector(to_unsigned(155, 8)),
			10658 => std_logic_vector(to_unsigned(102, 8)),
			10659 => std_logic_vector(to_unsigned(4, 8)),
			10660 => std_logic_vector(to_unsigned(84, 8)),
			10661 => std_logic_vector(to_unsigned(33, 8)),
			10662 => std_logic_vector(to_unsigned(213, 8)),
			10663 => std_logic_vector(to_unsigned(110, 8)),
			10664 => std_logic_vector(to_unsigned(100, 8)),
			10665 => std_logic_vector(to_unsigned(110, 8)),
			10666 => std_logic_vector(to_unsigned(83, 8)),
			10667 => std_logic_vector(to_unsigned(152, 8)),
			10668 => std_logic_vector(to_unsigned(40, 8)),
			10669 => std_logic_vector(to_unsigned(131, 8)),
			10670 => std_logic_vector(to_unsigned(16, 8)),
			10671 => std_logic_vector(to_unsigned(151, 8)),
			10672 => std_logic_vector(to_unsigned(187, 8)),
			10673 => std_logic_vector(to_unsigned(187, 8)),
			10674 => std_logic_vector(to_unsigned(183, 8)),
			10675 => std_logic_vector(to_unsigned(33, 8)),
			10676 => std_logic_vector(to_unsigned(242, 8)),
			10677 => std_logic_vector(to_unsigned(0, 8)),
			10678 => std_logic_vector(to_unsigned(76, 8)),
			10679 => std_logic_vector(to_unsigned(222, 8)),
			10680 => std_logic_vector(to_unsigned(147, 8)),
			10681 => std_logic_vector(to_unsigned(51, 8)),
			10682 => std_logic_vector(to_unsigned(149, 8)),
			10683 => std_logic_vector(to_unsigned(95, 8)),
			10684 => std_logic_vector(to_unsigned(77, 8)),
			10685 => std_logic_vector(to_unsigned(161, 8)),
			10686 => std_logic_vector(to_unsigned(10, 8)),
			10687 => std_logic_vector(to_unsigned(58, 8)),
			10688 => std_logic_vector(to_unsigned(16, 8)),
			10689 => std_logic_vector(to_unsigned(121, 8)),
			10690 => std_logic_vector(to_unsigned(68, 8)),
			10691 => std_logic_vector(to_unsigned(83, 8)),
			10692 => std_logic_vector(to_unsigned(154, 8)),
			10693 => std_logic_vector(to_unsigned(223, 8)),
			10694 => std_logic_vector(to_unsigned(62, 8)),
			10695 => std_logic_vector(to_unsigned(123, 8)),
			10696 => std_logic_vector(to_unsigned(127, 8)),
			10697 => std_logic_vector(to_unsigned(214, 8)),
			10698 => std_logic_vector(to_unsigned(102, 8)),
			10699 => std_logic_vector(to_unsigned(79, 8)),
			10700 => std_logic_vector(to_unsigned(195, 8)),
			10701 => std_logic_vector(to_unsigned(135, 8)),
			10702 => std_logic_vector(to_unsigned(49, 8)),
			10703 => std_logic_vector(to_unsigned(51, 8)),
			10704 => std_logic_vector(to_unsigned(189, 8)),
			10705 => std_logic_vector(to_unsigned(253, 8)),
			10706 => std_logic_vector(to_unsigned(122, 8)),
			10707 => std_logic_vector(to_unsigned(33, 8)),
			10708 => std_logic_vector(to_unsigned(45, 8)),
			10709 => std_logic_vector(to_unsigned(28, 8)),
			10710 => std_logic_vector(to_unsigned(170, 8)),
			10711 => std_logic_vector(to_unsigned(20, 8)),
			10712 => std_logic_vector(to_unsigned(229, 8)),
			10713 => std_logic_vector(to_unsigned(56, 8)),
			10714 => std_logic_vector(to_unsigned(30, 8)),
			10715 => std_logic_vector(to_unsigned(182, 8)),
			10716 => std_logic_vector(to_unsigned(180, 8)),
			10717 => std_logic_vector(to_unsigned(15, 8)),
			10718 => std_logic_vector(to_unsigned(189, 8)),
			10719 => std_logic_vector(to_unsigned(213, 8)),
			10720 => std_logic_vector(to_unsigned(199, 8)),
			10721 => std_logic_vector(to_unsigned(23, 8)),
			10722 => std_logic_vector(to_unsigned(184, 8)),
			10723 => std_logic_vector(to_unsigned(61, 8)),
			10724 => std_logic_vector(to_unsigned(208, 8)),
			10725 => std_logic_vector(to_unsigned(69, 8)),
			10726 => std_logic_vector(to_unsigned(26, 8)),
			10727 => std_logic_vector(to_unsigned(159, 8)),
			10728 => std_logic_vector(to_unsigned(142, 8)),
			10729 => std_logic_vector(to_unsigned(232, 8)),
			10730 => std_logic_vector(to_unsigned(120, 8)),
			10731 => std_logic_vector(to_unsigned(169, 8)),
			10732 => std_logic_vector(to_unsigned(33, 8)),
			10733 => std_logic_vector(to_unsigned(60, 8)),
			10734 => std_logic_vector(to_unsigned(213, 8)),
			10735 => std_logic_vector(to_unsigned(248, 8)),
			10736 => std_logic_vector(to_unsigned(158, 8)),
			10737 => std_logic_vector(to_unsigned(210, 8)),
			10738 => std_logic_vector(to_unsigned(98, 8)),
			10739 => std_logic_vector(to_unsigned(41, 8)),
			10740 => std_logic_vector(to_unsigned(37, 8)),
			10741 => std_logic_vector(to_unsigned(243, 8)),
			10742 => std_logic_vector(to_unsigned(1, 8)),
			10743 => std_logic_vector(to_unsigned(194, 8)),
			10744 => std_logic_vector(to_unsigned(19, 8)),
			10745 => std_logic_vector(to_unsigned(94, 8)),
			10746 => std_logic_vector(to_unsigned(90, 8)),
			10747 => std_logic_vector(to_unsigned(33, 8)),
			10748 => std_logic_vector(to_unsigned(234, 8)),
			10749 => std_logic_vector(to_unsigned(24, 8)),
			10750 => std_logic_vector(to_unsigned(199, 8)),
			10751 => std_logic_vector(to_unsigned(45, 8)),
			10752 => std_logic_vector(to_unsigned(78, 8)),
			10753 => std_logic_vector(to_unsigned(246, 8)),
			10754 => std_logic_vector(to_unsigned(104, 8)),
			10755 => std_logic_vector(to_unsigned(92, 8)),
			10756 => std_logic_vector(to_unsigned(64, 8)),
			10757 => std_logic_vector(to_unsigned(255, 8)),
			10758 => std_logic_vector(to_unsigned(233, 8)),
			10759 => std_logic_vector(to_unsigned(246, 8)),
			10760 => std_logic_vector(to_unsigned(248, 8)),
			10761 => std_logic_vector(to_unsigned(125, 8)),
			10762 => std_logic_vector(to_unsigned(46, 8)),
			10763 => std_logic_vector(to_unsigned(178, 8)),
			10764 => std_logic_vector(to_unsigned(87, 8)),
			10765 => std_logic_vector(to_unsigned(86, 8)),
			10766 => std_logic_vector(to_unsigned(147, 8)),
			10767 => std_logic_vector(to_unsigned(45, 8)),
			10768 => std_logic_vector(to_unsigned(72, 8)),
			10769 => std_logic_vector(to_unsigned(58, 8)),
			10770 => std_logic_vector(to_unsigned(8, 8)),
			10771 => std_logic_vector(to_unsigned(9, 8)),
			10772 => std_logic_vector(to_unsigned(171, 8)),
			10773 => std_logic_vector(to_unsigned(202, 8)),
			10774 => std_logic_vector(to_unsigned(5, 8)),
			10775 => std_logic_vector(to_unsigned(65, 8)),
			10776 => std_logic_vector(to_unsigned(128, 8)),
			10777 => std_logic_vector(to_unsigned(75, 8)),
			10778 => std_logic_vector(to_unsigned(67, 8)),
			10779 => std_logic_vector(to_unsigned(65, 8)),
			10780 => std_logic_vector(to_unsigned(245, 8)),
			10781 => std_logic_vector(to_unsigned(91, 8)),
			10782 => std_logic_vector(to_unsigned(1, 8)),
			10783 => std_logic_vector(to_unsigned(112, 8)),
			10784 => std_logic_vector(to_unsigned(123, 8)),
			10785 => std_logic_vector(to_unsigned(76, 8)),
			10786 => std_logic_vector(to_unsigned(168, 8)),
			10787 => std_logic_vector(to_unsigned(215, 8)),
			10788 => std_logic_vector(to_unsigned(17, 8)),
			10789 => std_logic_vector(to_unsigned(210, 8)),
			10790 => std_logic_vector(to_unsigned(247, 8)),
			10791 => std_logic_vector(to_unsigned(162, 8)),
			10792 => std_logic_vector(to_unsigned(238, 8)),
			10793 => std_logic_vector(to_unsigned(17, 8)),
			10794 => std_logic_vector(to_unsigned(48, 8)),
			10795 => std_logic_vector(to_unsigned(221, 8)),
			10796 => std_logic_vector(to_unsigned(17, 8)),
			10797 => std_logic_vector(to_unsigned(234, 8)),
			10798 => std_logic_vector(to_unsigned(192, 8)),
			10799 => std_logic_vector(to_unsigned(166, 8)),
			10800 => std_logic_vector(to_unsigned(138, 8)),
			10801 => std_logic_vector(to_unsigned(194, 8)),
			10802 => std_logic_vector(to_unsigned(193, 8)),
			10803 => std_logic_vector(to_unsigned(156, 8)),
			10804 => std_logic_vector(to_unsigned(108, 8)),
			10805 => std_logic_vector(to_unsigned(80, 8)),
			10806 => std_logic_vector(to_unsigned(10, 8)),
			10807 => std_logic_vector(to_unsigned(45, 8)),
			10808 => std_logic_vector(to_unsigned(0, 8)),
			10809 => std_logic_vector(to_unsigned(197, 8)),
			10810 => std_logic_vector(to_unsigned(53, 8)),
			10811 => std_logic_vector(to_unsigned(134, 8)),
			10812 => std_logic_vector(to_unsigned(96, 8)),
			10813 => std_logic_vector(to_unsigned(83, 8)),
			10814 => std_logic_vector(to_unsigned(118, 8)),
			10815 => std_logic_vector(to_unsigned(68, 8)),
			10816 => std_logic_vector(to_unsigned(129, 8)),
			10817 => std_logic_vector(to_unsigned(140, 8)),
			10818 => std_logic_vector(to_unsigned(161, 8)),
			10819 => std_logic_vector(to_unsigned(68, 8)),
			10820 => std_logic_vector(to_unsigned(41, 8)),
			10821 => std_logic_vector(to_unsigned(194, 8)),
			10822 => std_logic_vector(to_unsigned(138, 8)),
			10823 => std_logic_vector(to_unsigned(62, 8)),
			10824 => std_logic_vector(to_unsigned(136, 8)),
			10825 => std_logic_vector(to_unsigned(20, 8)),
			10826 => std_logic_vector(to_unsigned(176, 8)),
			10827 => std_logic_vector(to_unsigned(74, 8)),
			10828 => std_logic_vector(to_unsigned(190, 8)),
			10829 => std_logic_vector(to_unsigned(41, 8)),
			10830 => std_logic_vector(to_unsigned(200, 8)),
			10831 => std_logic_vector(to_unsigned(144, 8)),
			10832 => std_logic_vector(to_unsigned(77, 8)),
			10833 => std_logic_vector(to_unsigned(100, 8)),
			10834 => std_logic_vector(to_unsigned(168, 8)),
			10835 => std_logic_vector(to_unsigned(122, 8)),
			10836 => std_logic_vector(to_unsigned(111, 8)),
			10837 => std_logic_vector(to_unsigned(166, 8)),
			10838 => std_logic_vector(to_unsigned(228, 8)),
			10839 => std_logic_vector(to_unsigned(252, 8)),
			10840 => std_logic_vector(to_unsigned(65, 8)),
			10841 => std_logic_vector(to_unsigned(173, 8)),
			10842 => std_logic_vector(to_unsigned(27, 8)),
			10843 => std_logic_vector(to_unsigned(11, 8)),
			10844 => std_logic_vector(to_unsigned(118, 8)),
			10845 => std_logic_vector(to_unsigned(203, 8)),
			10846 => std_logic_vector(to_unsigned(9, 8)),
			10847 => std_logic_vector(to_unsigned(85, 8)),
			10848 => std_logic_vector(to_unsigned(252, 8)),
			10849 => std_logic_vector(to_unsigned(38, 8)),
			10850 => std_logic_vector(to_unsigned(42, 8)),
			10851 => std_logic_vector(to_unsigned(209, 8)),
			10852 => std_logic_vector(to_unsigned(84, 8)),
			10853 => std_logic_vector(to_unsigned(132, 8)),
			10854 => std_logic_vector(to_unsigned(71, 8)),
			10855 => std_logic_vector(to_unsigned(197, 8)),
			10856 => std_logic_vector(to_unsigned(110, 8)),
			10857 => std_logic_vector(to_unsigned(2, 8)),
			10858 => std_logic_vector(to_unsigned(93, 8)),
			10859 => std_logic_vector(to_unsigned(233, 8)),
			10860 => std_logic_vector(to_unsigned(1, 8)),
			10861 => std_logic_vector(to_unsigned(6, 8)),
			10862 => std_logic_vector(to_unsigned(101, 8)),
			10863 => std_logic_vector(to_unsigned(92, 8)),
			10864 => std_logic_vector(to_unsigned(197, 8)),
			10865 => std_logic_vector(to_unsigned(230, 8)),
			10866 => std_logic_vector(to_unsigned(170, 8)),
			10867 => std_logic_vector(to_unsigned(88, 8)),
			10868 => std_logic_vector(to_unsigned(147, 8)),
			10869 => std_logic_vector(to_unsigned(101, 8)),
			10870 => std_logic_vector(to_unsigned(131, 8)),
			10871 => std_logic_vector(to_unsigned(59, 8)),
			10872 => std_logic_vector(to_unsigned(31, 8)),
			10873 => std_logic_vector(to_unsigned(133, 8)),
			10874 => std_logic_vector(to_unsigned(98, 8)),
			10875 => std_logic_vector(to_unsigned(113, 8)),
			10876 => std_logic_vector(to_unsigned(69, 8)),
			10877 => std_logic_vector(to_unsigned(197, 8)),
			10878 => std_logic_vector(to_unsigned(21, 8)),
			10879 => std_logic_vector(to_unsigned(163, 8)),
			10880 => std_logic_vector(to_unsigned(224, 8)),
			10881 => std_logic_vector(to_unsigned(25, 8)),
			10882 => std_logic_vector(to_unsigned(42, 8)),
			10883 => std_logic_vector(to_unsigned(47, 8)),
			10884 => std_logic_vector(to_unsigned(4, 8)),
			10885 => std_logic_vector(to_unsigned(29, 8)),
			10886 => std_logic_vector(to_unsigned(227, 8)),
			10887 => std_logic_vector(to_unsigned(81, 8)),
			10888 => std_logic_vector(to_unsigned(114, 8)),
			10889 => std_logic_vector(to_unsigned(156, 8)),
			10890 => std_logic_vector(to_unsigned(255, 8)),
			10891 => std_logic_vector(to_unsigned(178, 8)),
			10892 => std_logic_vector(to_unsigned(246, 8)),
			10893 => std_logic_vector(to_unsigned(19, 8)),
			10894 => std_logic_vector(to_unsigned(246, 8)),
			10895 => std_logic_vector(to_unsigned(172, 8)),
			10896 => std_logic_vector(to_unsigned(63, 8)),
			10897 => std_logic_vector(to_unsigned(8, 8)),
			10898 => std_logic_vector(to_unsigned(5, 8)),
			10899 => std_logic_vector(to_unsigned(3, 8)),
			10900 => std_logic_vector(to_unsigned(9, 8)),
			10901 => std_logic_vector(to_unsigned(134, 8)),
			10902 => std_logic_vector(to_unsigned(62, 8)),
			10903 => std_logic_vector(to_unsigned(139, 8)),
			10904 => std_logic_vector(to_unsigned(240, 8)),
			10905 => std_logic_vector(to_unsigned(136, 8)),
			10906 => std_logic_vector(to_unsigned(186, 8)),
			10907 => std_logic_vector(to_unsigned(81, 8)),
			10908 => std_logic_vector(to_unsigned(44, 8)),
			10909 => std_logic_vector(to_unsigned(85, 8)),
			10910 => std_logic_vector(to_unsigned(224, 8)),
			10911 => std_logic_vector(to_unsigned(246, 8)),
			10912 => std_logic_vector(to_unsigned(33, 8)),
			10913 => std_logic_vector(to_unsigned(194, 8)),
			10914 => std_logic_vector(to_unsigned(147, 8)),
			10915 => std_logic_vector(to_unsigned(194, 8)),
			10916 => std_logic_vector(to_unsigned(43, 8)),
			10917 => std_logic_vector(to_unsigned(3, 8)),
			10918 => std_logic_vector(to_unsigned(48, 8)),
			10919 => std_logic_vector(to_unsigned(239, 8)),
			10920 => std_logic_vector(to_unsigned(222, 8)),
			10921 => std_logic_vector(to_unsigned(245, 8)),
			10922 => std_logic_vector(to_unsigned(163, 8)),
			10923 => std_logic_vector(to_unsigned(77, 8)),
			10924 => std_logic_vector(to_unsigned(251, 8)),
			10925 => std_logic_vector(to_unsigned(173, 8)),
			10926 => std_logic_vector(to_unsigned(238, 8)),
			10927 => std_logic_vector(to_unsigned(197, 8)),
			10928 => std_logic_vector(to_unsigned(170, 8)),
			10929 => std_logic_vector(to_unsigned(164, 8)),
			10930 => std_logic_vector(to_unsigned(37, 8)),
			10931 => std_logic_vector(to_unsigned(162, 8)),
			10932 => std_logic_vector(to_unsigned(13, 8)),
			10933 => std_logic_vector(to_unsigned(16, 8)),
			10934 => std_logic_vector(to_unsigned(34, 8)),
			10935 => std_logic_vector(to_unsigned(108, 8)),
			10936 => std_logic_vector(to_unsigned(146, 8)),
			10937 => std_logic_vector(to_unsigned(123, 8)),
			10938 => std_logic_vector(to_unsigned(218, 8)),
			10939 => std_logic_vector(to_unsigned(32, 8)),
			10940 => std_logic_vector(to_unsigned(100, 8)),
			10941 => std_logic_vector(to_unsigned(73, 8)),
			10942 => std_logic_vector(to_unsigned(58, 8)),
			10943 => std_logic_vector(to_unsigned(182, 8)),
			10944 => std_logic_vector(to_unsigned(132, 8)),
			10945 => std_logic_vector(to_unsigned(50, 8)),
			10946 => std_logic_vector(to_unsigned(30, 8)),
			10947 => std_logic_vector(to_unsigned(215, 8)),
			10948 => std_logic_vector(to_unsigned(32, 8)),
			10949 => std_logic_vector(to_unsigned(95, 8)),
			10950 => std_logic_vector(to_unsigned(237, 8)),
			10951 => std_logic_vector(to_unsigned(130, 8)),
			10952 => std_logic_vector(to_unsigned(237, 8)),
			10953 => std_logic_vector(to_unsigned(234, 8)),
			10954 => std_logic_vector(to_unsigned(137, 8)),
			10955 => std_logic_vector(to_unsigned(130, 8)),
			10956 => std_logic_vector(to_unsigned(68, 8)),
			10957 => std_logic_vector(to_unsigned(126, 8)),
			10958 => std_logic_vector(to_unsigned(112, 8)),
			10959 => std_logic_vector(to_unsigned(239, 8)),
			10960 => std_logic_vector(to_unsigned(97, 8)),
			10961 => std_logic_vector(to_unsigned(61, 8)),
			10962 => std_logic_vector(to_unsigned(153, 8)),
			10963 => std_logic_vector(to_unsigned(147, 8)),
			10964 => std_logic_vector(to_unsigned(30, 8)),
			10965 => std_logic_vector(to_unsigned(215, 8)),
			10966 => std_logic_vector(to_unsigned(185, 8)),
			10967 => std_logic_vector(to_unsigned(177, 8)),
			10968 => std_logic_vector(to_unsigned(182, 8)),
			10969 => std_logic_vector(to_unsigned(91, 8)),
			10970 => std_logic_vector(to_unsigned(139, 8)),
			10971 => std_logic_vector(to_unsigned(172, 8)),
			10972 => std_logic_vector(to_unsigned(52, 8)),
			10973 => std_logic_vector(to_unsigned(103, 8)),
			10974 => std_logic_vector(to_unsigned(77, 8)),
			10975 => std_logic_vector(to_unsigned(150, 8)),
			10976 => std_logic_vector(to_unsigned(95, 8)),
			10977 => std_logic_vector(to_unsigned(182, 8)),
			10978 => std_logic_vector(to_unsigned(214, 8)),
			10979 => std_logic_vector(to_unsigned(187, 8)),
			10980 => std_logic_vector(to_unsigned(247, 8)),
			10981 => std_logic_vector(to_unsigned(164, 8)),
			10982 => std_logic_vector(to_unsigned(184, 8)),
			10983 => std_logic_vector(to_unsigned(184, 8)),
			10984 => std_logic_vector(to_unsigned(166, 8)),
			10985 => std_logic_vector(to_unsigned(184, 8)),
			10986 => std_logic_vector(to_unsigned(112, 8)),
			10987 => std_logic_vector(to_unsigned(77, 8)),
			10988 => std_logic_vector(to_unsigned(122, 8)),
			10989 => std_logic_vector(to_unsigned(71, 8)),
			10990 => std_logic_vector(to_unsigned(141, 8)),
			10991 => std_logic_vector(to_unsigned(207, 8)),
			10992 => std_logic_vector(to_unsigned(45, 8)),
			10993 => std_logic_vector(to_unsigned(9, 8)),
			10994 => std_logic_vector(to_unsigned(201, 8)),
			10995 => std_logic_vector(to_unsigned(189, 8)),
			10996 => std_logic_vector(to_unsigned(121, 8)),
			10997 => std_logic_vector(to_unsigned(242, 8)),
			10998 => std_logic_vector(to_unsigned(104, 8)),
			10999 => std_logic_vector(to_unsigned(210, 8)),
			11000 => std_logic_vector(to_unsigned(85, 8)),
			11001 => std_logic_vector(to_unsigned(252, 8)),
			11002 => std_logic_vector(to_unsigned(217, 8)),
			11003 => std_logic_vector(to_unsigned(40, 8)),
			11004 => std_logic_vector(to_unsigned(250, 8)),
			11005 => std_logic_vector(to_unsigned(59, 8)),
			11006 => std_logic_vector(to_unsigned(183, 8)),
			11007 => std_logic_vector(to_unsigned(57, 8)),
			11008 => std_logic_vector(to_unsigned(151, 8)),
			11009 => std_logic_vector(to_unsigned(230, 8)),
			11010 => std_logic_vector(to_unsigned(7, 8)),
			11011 => std_logic_vector(to_unsigned(233, 8)),
			11012 => std_logic_vector(to_unsigned(227, 8)),
			11013 => std_logic_vector(to_unsigned(35, 8)),
			11014 => std_logic_vector(to_unsigned(90, 8)),
			11015 => std_logic_vector(to_unsigned(227, 8)),
			11016 => std_logic_vector(to_unsigned(145, 8)),
			11017 => std_logic_vector(to_unsigned(72, 8)),
			11018 => std_logic_vector(to_unsigned(36, 8)),
			11019 => std_logic_vector(to_unsigned(169, 8)),
			11020 => std_logic_vector(to_unsigned(57, 8)),
			11021 => std_logic_vector(to_unsigned(192, 8)),
			11022 => std_logic_vector(to_unsigned(18, 8)),
			11023 => std_logic_vector(to_unsigned(121, 8)),
			11024 => std_logic_vector(to_unsigned(28, 8)),
			11025 => std_logic_vector(to_unsigned(122, 8)),
			11026 => std_logic_vector(to_unsigned(216, 8)),
			11027 => std_logic_vector(to_unsigned(103, 8)),
			11028 => std_logic_vector(to_unsigned(221, 8)),
			11029 => std_logic_vector(to_unsigned(222, 8)),
			11030 => std_logic_vector(to_unsigned(197, 8)),
			11031 => std_logic_vector(to_unsigned(82, 8)),
			11032 => std_logic_vector(to_unsigned(218, 8)),
			11033 => std_logic_vector(to_unsigned(151, 8)),
			11034 => std_logic_vector(to_unsigned(141, 8)),
			11035 => std_logic_vector(to_unsigned(220, 8)),
			11036 => std_logic_vector(to_unsigned(240, 8)),
			11037 => std_logic_vector(to_unsigned(244, 8)),
			11038 => std_logic_vector(to_unsigned(177, 8)),
			11039 => std_logic_vector(to_unsigned(32, 8)),
			11040 => std_logic_vector(to_unsigned(117, 8)),
			11041 => std_logic_vector(to_unsigned(238, 8)),
			11042 => std_logic_vector(to_unsigned(204, 8)),
			11043 => std_logic_vector(to_unsigned(154, 8)),
			11044 => std_logic_vector(to_unsigned(231, 8)),
			11045 => std_logic_vector(to_unsigned(64, 8)),
			11046 => std_logic_vector(to_unsigned(6, 8)),
			11047 => std_logic_vector(to_unsigned(65, 8)),
			11048 => std_logic_vector(to_unsigned(78, 8)),
			11049 => std_logic_vector(to_unsigned(7, 8)),
			11050 => std_logic_vector(to_unsigned(175, 8)),
			11051 => std_logic_vector(to_unsigned(108, 8)),
			11052 => std_logic_vector(to_unsigned(125, 8)),
			11053 => std_logic_vector(to_unsigned(14, 8)),
			11054 => std_logic_vector(to_unsigned(118, 8)),
			11055 => std_logic_vector(to_unsigned(111, 8)),
			11056 => std_logic_vector(to_unsigned(204, 8)),
			11057 => std_logic_vector(to_unsigned(59, 8)),
			11058 => std_logic_vector(to_unsigned(7, 8)),
			11059 => std_logic_vector(to_unsigned(255, 8)),
			11060 => std_logic_vector(to_unsigned(158, 8)),
			11061 => std_logic_vector(to_unsigned(140, 8)),
			11062 => std_logic_vector(to_unsigned(220, 8)),
			11063 => std_logic_vector(to_unsigned(207, 8)),
			11064 => std_logic_vector(to_unsigned(73, 8)),
			11065 => std_logic_vector(to_unsigned(43, 8)),
			11066 => std_logic_vector(to_unsigned(225, 8)),
			11067 => std_logic_vector(to_unsigned(249, 8)),
			11068 => std_logic_vector(to_unsigned(169, 8)),
			11069 => std_logic_vector(to_unsigned(0, 8)),
			11070 => std_logic_vector(to_unsigned(151, 8)),
			11071 => std_logic_vector(to_unsigned(78, 8)),
			11072 => std_logic_vector(to_unsigned(23, 8)),
			11073 => std_logic_vector(to_unsigned(197, 8)),
			11074 => std_logic_vector(to_unsigned(65, 8)),
			11075 => std_logic_vector(to_unsigned(41, 8)),
			11076 => std_logic_vector(to_unsigned(242, 8)),
			11077 => std_logic_vector(to_unsigned(206, 8)),
			11078 => std_logic_vector(to_unsigned(192, 8)),
			11079 => std_logic_vector(to_unsigned(94, 8)),
			11080 => std_logic_vector(to_unsigned(39, 8)),
			11081 => std_logic_vector(to_unsigned(203, 8)),
			11082 => std_logic_vector(to_unsigned(2, 8)),
			11083 => std_logic_vector(to_unsigned(213, 8)),
			11084 => std_logic_vector(to_unsigned(124, 8)),
			11085 => std_logic_vector(to_unsigned(139, 8)),
			11086 => std_logic_vector(to_unsigned(87, 8)),
			11087 => std_logic_vector(to_unsigned(128, 8)),
			11088 => std_logic_vector(to_unsigned(176, 8)),
			11089 => std_logic_vector(to_unsigned(178, 8)),
			11090 => std_logic_vector(to_unsigned(239, 8)),
			11091 => std_logic_vector(to_unsigned(147, 8)),
			11092 => std_logic_vector(to_unsigned(136, 8)),
			11093 => std_logic_vector(to_unsigned(116, 8)),
			11094 => std_logic_vector(to_unsigned(120, 8)),
			11095 => std_logic_vector(to_unsigned(15, 8)),
			11096 => std_logic_vector(to_unsigned(100, 8)),
			11097 => std_logic_vector(to_unsigned(111, 8)),
			11098 => std_logic_vector(to_unsigned(179, 8)),
			11099 => std_logic_vector(to_unsigned(251, 8)),
			11100 => std_logic_vector(to_unsigned(234, 8)),
			11101 => std_logic_vector(to_unsigned(59, 8)),
			11102 => std_logic_vector(to_unsigned(46, 8)),
			11103 => std_logic_vector(to_unsigned(96, 8)),
			11104 => std_logic_vector(to_unsigned(33, 8)),
			11105 => std_logic_vector(to_unsigned(3, 8)),
			11106 => std_logic_vector(to_unsigned(179, 8)),
			11107 => std_logic_vector(to_unsigned(41, 8)),
			11108 => std_logic_vector(to_unsigned(131, 8)),
			11109 => std_logic_vector(to_unsigned(14, 8)),
			11110 => std_logic_vector(to_unsigned(20, 8)),
			11111 => std_logic_vector(to_unsigned(251, 8)),
			11112 => std_logic_vector(to_unsigned(131, 8)),
			11113 => std_logic_vector(to_unsigned(14, 8)),
			11114 => std_logic_vector(to_unsigned(116, 8)),
			11115 => std_logic_vector(to_unsigned(232, 8)),
			11116 => std_logic_vector(to_unsigned(94, 8)),
			11117 => std_logic_vector(to_unsigned(14, 8)),
			11118 => std_logic_vector(to_unsigned(71, 8)),
			11119 => std_logic_vector(to_unsigned(214, 8)),
			11120 => std_logic_vector(to_unsigned(106, 8)),
			11121 => std_logic_vector(to_unsigned(200, 8)),
			11122 => std_logic_vector(to_unsigned(204, 8)),
			11123 => std_logic_vector(to_unsigned(93, 8)),
			11124 => std_logic_vector(to_unsigned(158, 8)),
			11125 => std_logic_vector(to_unsigned(53, 8)),
			11126 => std_logic_vector(to_unsigned(241, 8)),
			11127 => std_logic_vector(to_unsigned(39, 8)),
			11128 => std_logic_vector(to_unsigned(36, 8)),
			11129 => std_logic_vector(to_unsigned(74, 8)),
			11130 => std_logic_vector(to_unsigned(132, 8)),
			11131 => std_logic_vector(to_unsigned(135, 8)),
			11132 => std_logic_vector(to_unsigned(163, 8)),
			11133 => std_logic_vector(to_unsigned(106, 8)),
			11134 => std_logic_vector(to_unsigned(33, 8)),
			11135 => std_logic_vector(to_unsigned(130, 8)),
			11136 => std_logic_vector(to_unsigned(164, 8)),
			11137 => std_logic_vector(to_unsigned(87, 8)),
			11138 => std_logic_vector(to_unsigned(198, 8)),
			11139 => std_logic_vector(to_unsigned(60, 8)),
			11140 => std_logic_vector(to_unsigned(82, 8)),
			11141 => std_logic_vector(to_unsigned(18, 8)),
			11142 => std_logic_vector(to_unsigned(231, 8)),
			11143 => std_logic_vector(to_unsigned(112, 8)),
			11144 => std_logic_vector(to_unsigned(43, 8)),
			11145 => std_logic_vector(to_unsigned(16, 8)),
			11146 => std_logic_vector(to_unsigned(185, 8)),
			11147 => std_logic_vector(to_unsigned(157, 8)),
			11148 => std_logic_vector(to_unsigned(40, 8)),
			11149 => std_logic_vector(to_unsigned(154, 8)),
			11150 => std_logic_vector(to_unsigned(174, 8)),
			11151 => std_logic_vector(to_unsigned(222, 8)),
			11152 => std_logic_vector(to_unsigned(196, 8)),
			11153 => std_logic_vector(to_unsigned(250, 8)),
			11154 => std_logic_vector(to_unsigned(159, 8)),
			11155 => std_logic_vector(to_unsigned(18, 8)),
			11156 => std_logic_vector(to_unsigned(30, 8)),
			11157 => std_logic_vector(to_unsigned(89, 8)),
			11158 => std_logic_vector(to_unsigned(36, 8)),
			11159 => std_logic_vector(to_unsigned(250, 8)),
			11160 => std_logic_vector(to_unsigned(164, 8)),
			11161 => std_logic_vector(to_unsigned(43, 8)),
			11162 => std_logic_vector(to_unsigned(96, 8)),
			11163 => std_logic_vector(to_unsigned(225, 8)),
			11164 => std_logic_vector(to_unsigned(240, 8)),
			11165 => std_logic_vector(to_unsigned(84, 8)),
			11166 => std_logic_vector(to_unsigned(205, 8)),
			11167 => std_logic_vector(to_unsigned(74, 8)),
			11168 => std_logic_vector(to_unsigned(50, 8)),
			11169 => std_logic_vector(to_unsigned(172, 8)),
			11170 => std_logic_vector(to_unsigned(68, 8)),
			11171 => std_logic_vector(to_unsigned(192, 8)),
			11172 => std_logic_vector(to_unsigned(224, 8)),
			11173 => std_logic_vector(to_unsigned(192, 8)),
			11174 => std_logic_vector(to_unsigned(1, 8)),
			11175 => std_logic_vector(to_unsigned(241, 8)),
			11176 => std_logic_vector(to_unsigned(189, 8)),
			11177 => std_logic_vector(to_unsigned(70, 8)),
			11178 => std_logic_vector(to_unsigned(222, 8)),
			11179 => std_logic_vector(to_unsigned(102, 8)),
			11180 => std_logic_vector(to_unsigned(147, 8)),
			11181 => std_logic_vector(to_unsigned(76, 8)),
			11182 => std_logic_vector(to_unsigned(145, 8)),
			11183 => std_logic_vector(to_unsigned(2, 8)),
			11184 => std_logic_vector(to_unsigned(186, 8)),
			11185 => std_logic_vector(to_unsigned(26, 8)),
			11186 => std_logic_vector(to_unsigned(135, 8)),
			11187 => std_logic_vector(to_unsigned(149, 8)),
			11188 => std_logic_vector(to_unsigned(232, 8)),
			11189 => std_logic_vector(to_unsigned(149, 8)),
			11190 => std_logic_vector(to_unsigned(44, 8)),
			11191 => std_logic_vector(to_unsigned(122, 8)),
			11192 => std_logic_vector(to_unsigned(61, 8)),
			11193 => std_logic_vector(to_unsigned(15, 8)),
			11194 => std_logic_vector(to_unsigned(228, 8)),
			11195 => std_logic_vector(to_unsigned(16, 8)),
			11196 => std_logic_vector(to_unsigned(96, 8)),
			11197 => std_logic_vector(to_unsigned(63, 8)),
			11198 => std_logic_vector(to_unsigned(208, 8)),
			11199 => std_logic_vector(to_unsigned(17, 8)),
			11200 => std_logic_vector(to_unsigned(194, 8)),
			11201 => std_logic_vector(to_unsigned(149, 8)),
			11202 => std_logic_vector(to_unsigned(204, 8)),
			11203 => std_logic_vector(to_unsigned(239, 8)),
			11204 => std_logic_vector(to_unsigned(133, 8)),
			11205 => std_logic_vector(to_unsigned(150, 8)),
			11206 => std_logic_vector(to_unsigned(3, 8)),
			11207 => std_logic_vector(to_unsigned(164, 8)),
			11208 => std_logic_vector(to_unsigned(8, 8)),
			11209 => std_logic_vector(to_unsigned(47, 8)),
			11210 => std_logic_vector(to_unsigned(197, 8)),
			11211 => std_logic_vector(to_unsigned(181, 8)),
			11212 => std_logic_vector(to_unsigned(36, 8)),
			11213 => std_logic_vector(to_unsigned(33, 8)),
			11214 => std_logic_vector(to_unsigned(255, 8)),
			11215 => std_logic_vector(to_unsigned(163, 8)),
			11216 => std_logic_vector(to_unsigned(31, 8)),
			11217 => std_logic_vector(to_unsigned(45, 8)),
			11218 => std_logic_vector(to_unsigned(240, 8)),
			11219 => std_logic_vector(to_unsigned(58, 8)),
			11220 => std_logic_vector(to_unsigned(232, 8)),
			11221 => std_logic_vector(to_unsigned(13, 8)),
			11222 => std_logic_vector(to_unsigned(40, 8)),
			11223 => std_logic_vector(to_unsigned(243, 8)),
			11224 => std_logic_vector(to_unsigned(168, 8)),
			11225 => std_logic_vector(to_unsigned(171, 8)),
			11226 => std_logic_vector(to_unsigned(32, 8)),
			11227 => std_logic_vector(to_unsigned(226, 8)),
			11228 => std_logic_vector(to_unsigned(243, 8)),
			11229 => std_logic_vector(to_unsigned(206, 8)),
			11230 => std_logic_vector(to_unsigned(0, 8)),
			11231 => std_logic_vector(to_unsigned(17, 8)),
			11232 => std_logic_vector(to_unsigned(167, 8)),
			11233 => std_logic_vector(to_unsigned(31, 8)),
			11234 => std_logic_vector(to_unsigned(10, 8)),
			11235 => std_logic_vector(to_unsigned(164, 8)),
			11236 => std_logic_vector(to_unsigned(213, 8)),
			11237 => std_logic_vector(to_unsigned(255, 8)),
			11238 => std_logic_vector(to_unsigned(50, 8)),
			11239 => std_logic_vector(to_unsigned(161, 8)),
			11240 => std_logic_vector(to_unsigned(93, 8)),
			11241 => std_logic_vector(to_unsigned(14, 8)),
			11242 => std_logic_vector(to_unsigned(48, 8)),
			11243 => std_logic_vector(to_unsigned(249, 8)),
			11244 => std_logic_vector(to_unsigned(212, 8)),
			11245 => std_logic_vector(to_unsigned(57, 8)),
			11246 => std_logic_vector(to_unsigned(171, 8)),
			11247 => std_logic_vector(to_unsigned(106, 8)),
			11248 => std_logic_vector(to_unsigned(14, 8)),
			11249 => std_logic_vector(to_unsigned(129, 8)),
			11250 => std_logic_vector(to_unsigned(183, 8)),
			11251 => std_logic_vector(to_unsigned(165, 8)),
			11252 => std_logic_vector(to_unsigned(100, 8)),
			11253 => std_logic_vector(to_unsigned(208, 8)),
			11254 => std_logic_vector(to_unsigned(244, 8)),
			11255 => std_logic_vector(to_unsigned(45, 8)),
			11256 => std_logic_vector(to_unsigned(96, 8)),
			11257 => std_logic_vector(to_unsigned(166, 8)),
			11258 => std_logic_vector(to_unsigned(120, 8)),
			11259 => std_logic_vector(to_unsigned(3, 8)),
			11260 => std_logic_vector(to_unsigned(29, 8)),
			11261 => std_logic_vector(to_unsigned(225, 8)),
			11262 => std_logic_vector(to_unsigned(251, 8)),
			11263 => std_logic_vector(to_unsigned(211, 8)),
			11264 => std_logic_vector(to_unsigned(253, 8)),
			11265 => std_logic_vector(to_unsigned(16, 8)),
			11266 => std_logic_vector(to_unsigned(92, 8)),
			11267 => std_logic_vector(to_unsigned(230, 8)),
			11268 => std_logic_vector(to_unsigned(198, 8)),
			11269 => std_logic_vector(to_unsigned(124, 8)),
			11270 => std_logic_vector(to_unsigned(149, 8)),
			11271 => std_logic_vector(to_unsigned(120, 8)),
			11272 => std_logic_vector(to_unsigned(86, 8)),
			11273 => std_logic_vector(to_unsigned(144, 8)),
			11274 => std_logic_vector(to_unsigned(17, 8)),
			11275 => std_logic_vector(to_unsigned(255, 8)),
			11276 => std_logic_vector(to_unsigned(106, 8)),
			11277 => std_logic_vector(to_unsigned(230, 8)),
			11278 => std_logic_vector(to_unsigned(22, 8)),
			11279 => std_logic_vector(to_unsigned(210, 8)),
			11280 => std_logic_vector(to_unsigned(80, 8)),
			11281 => std_logic_vector(to_unsigned(91, 8)),
			11282 => std_logic_vector(to_unsigned(243, 8)),
			11283 => std_logic_vector(to_unsigned(126, 8)),
			11284 => std_logic_vector(to_unsigned(161, 8)),
			11285 => std_logic_vector(to_unsigned(181, 8)),
			11286 => std_logic_vector(to_unsigned(246, 8)),
			11287 => std_logic_vector(to_unsigned(26, 8)),
			11288 => std_logic_vector(to_unsigned(240, 8)),
			11289 => std_logic_vector(to_unsigned(235, 8)),
			11290 => std_logic_vector(to_unsigned(178, 8)),
			11291 => std_logic_vector(to_unsigned(19, 8)),
			11292 => std_logic_vector(to_unsigned(113, 8)),
			11293 => std_logic_vector(to_unsigned(152, 8)),
			11294 => std_logic_vector(to_unsigned(86, 8)),
			11295 => std_logic_vector(to_unsigned(127, 8)),
			11296 => std_logic_vector(to_unsigned(224, 8)),
			11297 => std_logic_vector(to_unsigned(44, 8)),
			11298 => std_logic_vector(to_unsigned(212, 8)),
			11299 => std_logic_vector(to_unsigned(187, 8)),
			11300 => std_logic_vector(to_unsigned(1, 8)),
			11301 => std_logic_vector(to_unsigned(241, 8)),
			11302 => std_logic_vector(to_unsigned(108, 8)),
			11303 => std_logic_vector(to_unsigned(35, 8)),
			11304 => std_logic_vector(to_unsigned(28, 8)),
			11305 => std_logic_vector(to_unsigned(8, 8)),
			11306 => std_logic_vector(to_unsigned(74, 8)),
			11307 => std_logic_vector(to_unsigned(32, 8)),
			11308 => std_logic_vector(to_unsigned(250, 8)),
			11309 => std_logic_vector(to_unsigned(174, 8)),
			11310 => std_logic_vector(to_unsigned(46, 8)),
			11311 => std_logic_vector(to_unsigned(119, 8)),
			11312 => std_logic_vector(to_unsigned(19, 8)),
			11313 => std_logic_vector(to_unsigned(67, 8)),
			11314 => std_logic_vector(to_unsigned(66, 8)),
			11315 => std_logic_vector(to_unsigned(247, 8)),
			11316 => std_logic_vector(to_unsigned(187, 8)),
			11317 => std_logic_vector(to_unsigned(130, 8)),
			11318 => std_logic_vector(to_unsigned(212, 8)),
			11319 => std_logic_vector(to_unsigned(13, 8)),
			11320 => std_logic_vector(to_unsigned(183, 8)),
			11321 => std_logic_vector(to_unsigned(69, 8)),
			11322 => std_logic_vector(to_unsigned(246, 8)),
			11323 => std_logic_vector(to_unsigned(216, 8)),
			11324 => std_logic_vector(to_unsigned(253, 8)),
			11325 => std_logic_vector(to_unsigned(172, 8)),
			11326 => std_logic_vector(to_unsigned(3, 8)),
			11327 => std_logic_vector(to_unsigned(158, 8)),
			11328 => std_logic_vector(to_unsigned(10, 8)),
			11329 => std_logic_vector(to_unsigned(60, 8)),
			11330 => std_logic_vector(to_unsigned(49, 8)),
			11331 => std_logic_vector(to_unsigned(165, 8)),
			11332 => std_logic_vector(to_unsigned(55, 8)),
			11333 => std_logic_vector(to_unsigned(150, 8)),
			11334 => std_logic_vector(to_unsigned(101, 8)),
			11335 => std_logic_vector(to_unsigned(70, 8)),
			11336 => std_logic_vector(to_unsigned(136, 8)),
			11337 => std_logic_vector(to_unsigned(70, 8)),
			11338 => std_logic_vector(to_unsigned(73, 8)),
			11339 => std_logic_vector(to_unsigned(153, 8)),
			11340 => std_logic_vector(to_unsigned(252, 8)),
			11341 => std_logic_vector(to_unsigned(123, 8)),
			11342 => std_logic_vector(to_unsigned(45, 8)),
			11343 => std_logic_vector(to_unsigned(235, 8)),
			11344 => std_logic_vector(to_unsigned(132, 8)),
			11345 => std_logic_vector(to_unsigned(181, 8)),
			11346 => std_logic_vector(to_unsigned(40, 8)),
			11347 => std_logic_vector(to_unsigned(143, 8)),
			11348 => std_logic_vector(to_unsigned(87, 8)),
			11349 => std_logic_vector(to_unsigned(109, 8)),
			11350 => std_logic_vector(to_unsigned(243, 8)),
			11351 => std_logic_vector(to_unsigned(87, 8)),
			11352 => std_logic_vector(to_unsigned(121, 8)),
			11353 => std_logic_vector(to_unsigned(251, 8)),
			11354 => std_logic_vector(to_unsigned(164, 8)),
			11355 => std_logic_vector(to_unsigned(156, 8)),
			11356 => std_logic_vector(to_unsigned(23, 8)),
			11357 => std_logic_vector(to_unsigned(59, 8)),
			11358 => std_logic_vector(to_unsigned(72, 8)),
			11359 => std_logic_vector(to_unsigned(106, 8)),
			11360 => std_logic_vector(to_unsigned(219, 8)),
			11361 => std_logic_vector(to_unsigned(3, 8)),
			11362 => std_logic_vector(to_unsigned(52, 8)),
			11363 => std_logic_vector(to_unsigned(166, 8)),
			11364 => std_logic_vector(to_unsigned(183, 8)),
			11365 => std_logic_vector(to_unsigned(214, 8)),
			11366 => std_logic_vector(to_unsigned(197, 8)),
			11367 => std_logic_vector(to_unsigned(227, 8)),
			11368 => std_logic_vector(to_unsigned(45, 8)),
			11369 => std_logic_vector(to_unsigned(216, 8)),
			11370 => std_logic_vector(to_unsigned(98, 8)),
			11371 => std_logic_vector(to_unsigned(193, 8)),
			11372 => std_logic_vector(to_unsigned(131, 8)),
			11373 => std_logic_vector(to_unsigned(18, 8)),
			11374 => std_logic_vector(to_unsigned(126, 8)),
			11375 => std_logic_vector(to_unsigned(242, 8)),
			11376 => std_logic_vector(to_unsigned(19, 8)),
			11377 => std_logic_vector(to_unsigned(27, 8)),
			11378 => std_logic_vector(to_unsigned(255, 8)),
			11379 => std_logic_vector(to_unsigned(103, 8)),
			11380 => std_logic_vector(to_unsigned(176, 8)),
			11381 => std_logic_vector(to_unsigned(163, 8)),
			11382 => std_logic_vector(to_unsigned(193, 8)),
			11383 => std_logic_vector(to_unsigned(125, 8)),
			11384 => std_logic_vector(to_unsigned(29, 8)),
			11385 => std_logic_vector(to_unsigned(204, 8)),
			11386 => std_logic_vector(to_unsigned(110, 8)),
			11387 => std_logic_vector(to_unsigned(242, 8)),
			11388 => std_logic_vector(to_unsigned(137, 8)),
			11389 => std_logic_vector(to_unsigned(171, 8)),
			11390 => std_logic_vector(to_unsigned(250, 8)),
			11391 => std_logic_vector(to_unsigned(176, 8)),
			11392 => std_logic_vector(to_unsigned(242, 8)),
			11393 => std_logic_vector(to_unsigned(133, 8)),
			11394 => std_logic_vector(to_unsigned(12, 8)),
			11395 => std_logic_vector(to_unsigned(63, 8)),
			11396 => std_logic_vector(to_unsigned(111, 8)),
			11397 => std_logic_vector(to_unsigned(191, 8)),
			11398 => std_logic_vector(to_unsigned(118, 8)),
			11399 => std_logic_vector(to_unsigned(73, 8)),
			11400 => std_logic_vector(to_unsigned(14, 8)),
			11401 => std_logic_vector(to_unsigned(77, 8)),
			11402 => std_logic_vector(to_unsigned(136, 8)),
			11403 => std_logic_vector(to_unsigned(141, 8)),
			11404 => std_logic_vector(to_unsigned(188, 8)),
			11405 => std_logic_vector(to_unsigned(219, 8)),
			11406 => std_logic_vector(to_unsigned(37, 8)),
			11407 => std_logic_vector(to_unsigned(100, 8)),
			11408 => std_logic_vector(to_unsigned(105, 8)),
			11409 => std_logic_vector(to_unsigned(236, 8)),
			11410 => std_logic_vector(to_unsigned(162, 8)),
			11411 => std_logic_vector(to_unsigned(142, 8)),
			11412 => std_logic_vector(to_unsigned(218, 8)),
			11413 => std_logic_vector(to_unsigned(159, 8)),
			11414 => std_logic_vector(to_unsigned(233, 8)),
			11415 => std_logic_vector(to_unsigned(208, 8)),
			11416 => std_logic_vector(to_unsigned(4, 8)),
			11417 => std_logic_vector(to_unsigned(190, 8)),
			11418 => std_logic_vector(to_unsigned(180, 8)),
			11419 => std_logic_vector(to_unsigned(180, 8)),
			11420 => std_logic_vector(to_unsigned(128, 8)),
			11421 => std_logic_vector(to_unsigned(57, 8)),
			11422 => std_logic_vector(to_unsigned(64, 8)),
			11423 => std_logic_vector(to_unsigned(157, 8)),
			11424 => std_logic_vector(to_unsigned(246, 8)),
			11425 => std_logic_vector(to_unsigned(38, 8)),
			11426 => std_logic_vector(to_unsigned(19, 8)),
			11427 => std_logic_vector(to_unsigned(199, 8)),
			11428 => std_logic_vector(to_unsigned(249, 8)),
			11429 => std_logic_vector(to_unsigned(15, 8)),
			11430 => std_logic_vector(to_unsigned(175, 8)),
			11431 => std_logic_vector(to_unsigned(215, 8)),
			11432 => std_logic_vector(to_unsigned(3, 8)),
			11433 => std_logic_vector(to_unsigned(98, 8)),
			11434 => std_logic_vector(to_unsigned(68, 8)),
			11435 => std_logic_vector(to_unsigned(247, 8)),
			11436 => std_logic_vector(to_unsigned(39, 8)),
			11437 => std_logic_vector(to_unsigned(139, 8)),
			11438 => std_logic_vector(to_unsigned(39, 8)),
			11439 => std_logic_vector(to_unsigned(161, 8)),
			11440 => std_logic_vector(to_unsigned(142, 8)),
			11441 => std_logic_vector(to_unsigned(149, 8)),
			11442 => std_logic_vector(to_unsigned(79, 8)),
			11443 => std_logic_vector(to_unsigned(121, 8)),
			11444 => std_logic_vector(to_unsigned(24, 8)),
			11445 => std_logic_vector(to_unsigned(102, 8)),
			11446 => std_logic_vector(to_unsigned(111, 8)),
			11447 => std_logic_vector(to_unsigned(2, 8)),
			11448 => std_logic_vector(to_unsigned(227, 8)),
			11449 => std_logic_vector(to_unsigned(39, 8)),
			11450 => std_logic_vector(to_unsigned(52, 8)),
			11451 => std_logic_vector(to_unsigned(77, 8)),
			11452 => std_logic_vector(to_unsigned(130, 8)),
			11453 => std_logic_vector(to_unsigned(12, 8)),
			11454 => std_logic_vector(to_unsigned(156, 8)),
			11455 => std_logic_vector(to_unsigned(205, 8)),
			11456 => std_logic_vector(to_unsigned(31, 8)),
			11457 => std_logic_vector(to_unsigned(126, 8)),
			11458 => std_logic_vector(to_unsigned(61, 8)),
			11459 => std_logic_vector(to_unsigned(155, 8)),
			11460 => std_logic_vector(to_unsigned(31, 8)),
			11461 => std_logic_vector(to_unsigned(238, 8)),
			11462 => std_logic_vector(to_unsigned(138, 8)),
			11463 => std_logic_vector(to_unsigned(104, 8)),
			11464 => std_logic_vector(to_unsigned(58, 8)),
			11465 => std_logic_vector(to_unsigned(81, 8)),
			11466 => std_logic_vector(to_unsigned(214, 8)),
			11467 => std_logic_vector(to_unsigned(56, 8)),
			11468 => std_logic_vector(to_unsigned(169, 8)),
			11469 => std_logic_vector(to_unsigned(207, 8)),
			11470 => std_logic_vector(to_unsigned(189, 8)),
			11471 => std_logic_vector(to_unsigned(228, 8)),
			11472 => std_logic_vector(to_unsigned(64, 8)),
			11473 => std_logic_vector(to_unsigned(148, 8)),
			11474 => std_logic_vector(to_unsigned(70, 8)),
			11475 => std_logic_vector(to_unsigned(104, 8)),
			11476 => std_logic_vector(to_unsigned(125, 8)),
			11477 => std_logic_vector(to_unsigned(250, 8)),
			11478 => std_logic_vector(to_unsigned(121, 8)),
			11479 => std_logic_vector(to_unsigned(102, 8)),
			11480 => std_logic_vector(to_unsigned(242, 8)),
			11481 => std_logic_vector(to_unsigned(195, 8)),
			11482 => std_logic_vector(to_unsigned(20, 8)),
			11483 => std_logic_vector(to_unsigned(68, 8)),
			11484 => std_logic_vector(to_unsigned(243, 8)),
			11485 => std_logic_vector(to_unsigned(252, 8)),
			11486 => std_logic_vector(to_unsigned(188, 8)),
			11487 => std_logic_vector(to_unsigned(244, 8)),
			11488 => std_logic_vector(to_unsigned(1, 8)),
			11489 => std_logic_vector(to_unsigned(133, 8)),
			11490 => std_logic_vector(to_unsigned(194, 8)),
			11491 => std_logic_vector(to_unsigned(56, 8)),
			11492 => std_logic_vector(to_unsigned(146, 8)),
			11493 => std_logic_vector(to_unsigned(98, 8)),
			11494 => std_logic_vector(to_unsigned(178, 8)),
			11495 => std_logic_vector(to_unsigned(109, 8)),
			11496 => std_logic_vector(to_unsigned(62, 8)),
			11497 => std_logic_vector(to_unsigned(185, 8)),
			11498 => std_logic_vector(to_unsigned(35, 8)),
			11499 => std_logic_vector(to_unsigned(121, 8)),
			11500 => std_logic_vector(to_unsigned(127, 8)),
			11501 => std_logic_vector(to_unsigned(9, 8)),
			11502 => std_logic_vector(to_unsigned(194, 8)),
			11503 => std_logic_vector(to_unsigned(129, 8)),
			11504 => std_logic_vector(to_unsigned(217, 8)),
			11505 => std_logic_vector(to_unsigned(82, 8)),
			11506 => std_logic_vector(to_unsigned(30, 8)),
			11507 => std_logic_vector(to_unsigned(175, 8)),
			11508 => std_logic_vector(to_unsigned(17, 8)),
			11509 => std_logic_vector(to_unsigned(42, 8)),
			11510 => std_logic_vector(to_unsigned(49, 8)),
			11511 => std_logic_vector(to_unsigned(245, 8)),
			11512 => std_logic_vector(to_unsigned(62, 8)),
			11513 => std_logic_vector(to_unsigned(155, 8)),
			11514 => std_logic_vector(to_unsigned(23, 8)),
			11515 => std_logic_vector(to_unsigned(51, 8)),
			11516 => std_logic_vector(to_unsigned(203, 8)),
			11517 => std_logic_vector(to_unsigned(233, 8)),
			11518 => std_logic_vector(to_unsigned(244, 8)),
			11519 => std_logic_vector(to_unsigned(233, 8)),
			11520 => std_logic_vector(to_unsigned(194, 8)),
			11521 => std_logic_vector(to_unsigned(174, 8)),
			11522 => std_logic_vector(to_unsigned(131, 8)),
			11523 => std_logic_vector(to_unsigned(155, 8)),
			11524 => std_logic_vector(to_unsigned(57, 8)),
			11525 => std_logic_vector(to_unsigned(158, 8)),
			11526 => std_logic_vector(to_unsigned(226, 8)),
			11527 => std_logic_vector(to_unsigned(151, 8)),
			11528 => std_logic_vector(to_unsigned(138, 8)),
			11529 => std_logic_vector(to_unsigned(53, 8)),
			11530 => std_logic_vector(to_unsigned(233, 8)),
			11531 => std_logic_vector(to_unsigned(64, 8)),
			11532 => std_logic_vector(to_unsigned(137, 8)),
			11533 => std_logic_vector(to_unsigned(176, 8)),
			11534 => std_logic_vector(to_unsigned(194, 8)),
			11535 => std_logic_vector(to_unsigned(124, 8)),
			11536 => std_logic_vector(to_unsigned(13, 8)),
			11537 => std_logic_vector(to_unsigned(70, 8)),
			11538 => std_logic_vector(to_unsigned(226, 8)),
			11539 => std_logic_vector(to_unsigned(139, 8)),
			11540 => std_logic_vector(to_unsigned(217, 8)),
			11541 => std_logic_vector(to_unsigned(174, 8)),
			11542 => std_logic_vector(to_unsigned(136, 8)),
			11543 => std_logic_vector(to_unsigned(212, 8)),
			11544 => std_logic_vector(to_unsigned(176, 8)),
			11545 => std_logic_vector(to_unsigned(235, 8)),
			11546 => std_logic_vector(to_unsigned(69, 8)),
			11547 => std_logic_vector(to_unsigned(87, 8)),
			11548 => std_logic_vector(to_unsigned(75, 8)),
			11549 => std_logic_vector(to_unsigned(192, 8)),
			11550 => std_logic_vector(to_unsigned(58, 8)),
			11551 => std_logic_vector(to_unsigned(100, 8)),
			11552 => std_logic_vector(to_unsigned(65, 8)),
			11553 => std_logic_vector(to_unsigned(113, 8)),
			11554 => std_logic_vector(to_unsigned(44, 8)),
			11555 => std_logic_vector(to_unsigned(112, 8)),
			11556 => std_logic_vector(to_unsigned(102, 8)),
			11557 => std_logic_vector(to_unsigned(95, 8)),
			11558 => std_logic_vector(to_unsigned(82, 8)),
			11559 => std_logic_vector(to_unsigned(137, 8)),
			11560 => std_logic_vector(to_unsigned(81, 8)),
			11561 => std_logic_vector(to_unsigned(158, 8)),
			11562 => std_logic_vector(to_unsigned(82, 8)),
			11563 => std_logic_vector(to_unsigned(2, 8)),
			11564 => std_logic_vector(to_unsigned(123, 8)),
			11565 => std_logic_vector(to_unsigned(178, 8)),
			11566 => std_logic_vector(to_unsigned(167, 8)),
			11567 => std_logic_vector(to_unsigned(172, 8)),
			11568 => std_logic_vector(to_unsigned(239, 8)),
			11569 => std_logic_vector(to_unsigned(24, 8)),
			11570 => std_logic_vector(to_unsigned(199, 8)),
			11571 => std_logic_vector(to_unsigned(15, 8)),
			11572 => std_logic_vector(to_unsigned(161, 8)),
			11573 => std_logic_vector(to_unsigned(222, 8)),
			11574 => std_logic_vector(to_unsigned(183, 8)),
			11575 => std_logic_vector(to_unsigned(19, 8)),
			11576 => std_logic_vector(to_unsigned(54, 8)),
			11577 => std_logic_vector(to_unsigned(254, 8)),
			11578 => std_logic_vector(to_unsigned(61, 8)),
			11579 => std_logic_vector(to_unsigned(233, 8)),
			11580 => std_logic_vector(to_unsigned(141, 8)),
			11581 => std_logic_vector(to_unsigned(47, 8)),
			11582 => std_logic_vector(to_unsigned(11, 8)),
			11583 => std_logic_vector(to_unsigned(170, 8)),
			11584 => std_logic_vector(to_unsigned(225, 8)),
			11585 => std_logic_vector(to_unsigned(1, 8)),
			11586 => std_logic_vector(to_unsigned(126, 8)),
			11587 => std_logic_vector(to_unsigned(135, 8)),
			11588 => std_logic_vector(to_unsigned(69, 8)),
			11589 => std_logic_vector(to_unsigned(83, 8)),
			11590 => std_logic_vector(to_unsigned(179, 8)),
			11591 => std_logic_vector(to_unsigned(147, 8)),
			11592 => std_logic_vector(to_unsigned(28, 8)),
			11593 => std_logic_vector(to_unsigned(98, 8)),
			11594 => std_logic_vector(to_unsigned(119, 8)),
			11595 => std_logic_vector(to_unsigned(108, 8)),
			11596 => std_logic_vector(to_unsigned(19, 8)),
			11597 => std_logic_vector(to_unsigned(188, 8)),
			11598 => std_logic_vector(to_unsigned(249, 8)),
			11599 => std_logic_vector(to_unsigned(69, 8)),
			11600 => std_logic_vector(to_unsigned(174, 8)),
			11601 => std_logic_vector(to_unsigned(86, 8)),
			11602 => std_logic_vector(to_unsigned(215, 8)),
			11603 => std_logic_vector(to_unsigned(25, 8)),
			11604 => std_logic_vector(to_unsigned(72, 8)),
			11605 => std_logic_vector(to_unsigned(199, 8)),
			11606 => std_logic_vector(to_unsigned(204, 8)),
			11607 => std_logic_vector(to_unsigned(123, 8)),
			11608 => std_logic_vector(to_unsigned(125, 8)),
			11609 => std_logic_vector(to_unsigned(1, 8)),
			11610 => std_logic_vector(to_unsigned(231, 8)),
			11611 => std_logic_vector(to_unsigned(116, 8)),
			11612 => std_logic_vector(to_unsigned(117, 8)),
			11613 => std_logic_vector(to_unsigned(1, 8)),
			11614 => std_logic_vector(to_unsigned(106, 8)),
			11615 => std_logic_vector(to_unsigned(229, 8)),
			11616 => std_logic_vector(to_unsigned(100, 8)),
			11617 => std_logic_vector(to_unsigned(192, 8)),
			11618 => std_logic_vector(to_unsigned(146, 8)),
			11619 => std_logic_vector(to_unsigned(253, 8)),
			11620 => std_logic_vector(to_unsigned(231, 8)),
			11621 => std_logic_vector(to_unsigned(115, 8)),
			11622 => std_logic_vector(to_unsigned(249, 8)),
			11623 => std_logic_vector(to_unsigned(142, 8)),
			11624 => std_logic_vector(to_unsigned(252, 8)),
			11625 => std_logic_vector(to_unsigned(104, 8)),
			11626 => std_logic_vector(to_unsigned(216, 8)),
			11627 => std_logic_vector(to_unsigned(108, 8)),
			11628 => std_logic_vector(to_unsigned(96, 8)),
			11629 => std_logic_vector(to_unsigned(39, 8)),
			11630 => std_logic_vector(to_unsigned(43, 8)),
			11631 => std_logic_vector(to_unsigned(58, 8)),
			11632 => std_logic_vector(to_unsigned(129, 8)),
			11633 => std_logic_vector(to_unsigned(73, 8)),
			11634 => std_logic_vector(to_unsigned(169, 8)),
			11635 => std_logic_vector(to_unsigned(55, 8)),
			11636 => std_logic_vector(to_unsigned(166, 8)),
			11637 => std_logic_vector(to_unsigned(21, 8)),
			11638 => std_logic_vector(to_unsigned(241, 8)),
			11639 => std_logic_vector(to_unsigned(118, 8)),
			11640 => std_logic_vector(to_unsigned(68, 8)),
			11641 => std_logic_vector(to_unsigned(134, 8)),
			others => (others => '0'));
component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;
begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;
MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end process;
test : process is
begin 
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;
	assert RAM(11642) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(11642))))  severity failure;
	assert RAM(11643) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(11643))))  severity failure;
	assert RAM(11644) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(11644))))  severity failure;
	assert RAM(11645) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(11645))))  severity failure;
	assert RAM(11646) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(11646))))  severity failure;
	assert RAM(11647) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(11647))))  severity failure;
	assert RAM(11648) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(11648))))  severity failure;
	assert RAM(11649) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(11649))))  severity failure;
	assert RAM(11650) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(11650))))  severity failure;
	assert RAM(11651) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(11651))))  severity failure;
	assert RAM(11652) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(11652))))  severity failure;
	assert RAM(11653) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(11653))))  severity failure;
	assert RAM(11654) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(11654))))  severity failure;
	assert RAM(11655) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(11655))))  severity failure;
	assert RAM(11656) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(11656))))  severity failure;
	assert RAM(11657) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(11657))))  severity failure;
	assert RAM(11658) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(11658))))  severity failure;
	assert RAM(11659) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(11659))))  severity failure;
	assert RAM(11660) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(11660))))  severity failure;
	assert RAM(11661) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(11661))))  severity failure;
	assert RAM(11662) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(11662))))  severity failure;
	assert RAM(11663) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(11663))))  severity failure;
	assert RAM(11664) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(11664))))  severity failure;
	assert RAM(11665) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(11665))))  severity failure;
	assert RAM(11666) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(11666))))  severity failure;
	assert RAM(11667) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(11667))))  severity failure;
	assert RAM(11668) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(11668))))  severity failure;
	assert RAM(11669) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(11669))))  severity failure;
	assert RAM(11670) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(11670))))  severity failure;
	assert RAM(11671) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(11671))))  severity failure;
	assert RAM(11672) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(11672))))  severity failure;
	assert RAM(11673) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(11673))))  severity failure;
	assert RAM(11674) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(11674))))  severity failure;
	assert RAM(11675) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(11675))))  severity failure;
	assert RAM(11676) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(11676))))  severity failure;
	assert RAM(11677) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(11677))))  severity failure;
	assert RAM(11678) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(11678))))  severity failure;
	assert RAM(11679) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(11679))))  severity failure;
	assert RAM(11680) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(11680))))  severity failure;
	assert RAM(11681) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(11681))))  severity failure;
	assert RAM(11682) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(11682))))  severity failure;
	assert RAM(11683) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(11683))))  severity failure;
	assert RAM(11684) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(11684))))  severity failure;
	assert RAM(11685) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(11685))))  severity failure;
	assert RAM(11686) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(11686))))  severity failure;
	assert RAM(11687) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(11687))))  severity failure;
	assert RAM(11688) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(11688))))  severity failure;
	assert RAM(11689) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(11689))))  severity failure;
	assert RAM(11690) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(11690))))  severity failure;
	assert RAM(11691) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(11691))))  severity failure;
	assert RAM(11692) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(11692))))  severity failure;
	assert RAM(11693) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(11693))))  severity failure;
	assert RAM(11694) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(11694))))  severity failure;
	assert RAM(11695) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(11695))))  severity failure;
	assert RAM(11696) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(11696))))  severity failure;
	assert RAM(11697) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(11697))))  severity failure;
	assert RAM(11698) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(11698))))  severity failure;
	assert RAM(11699) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(11699))))  severity failure;
	assert RAM(11700) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(11700))))  severity failure;
	assert RAM(11701) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(11701))))  severity failure;
	assert RAM(11702) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(11702))))  severity failure;
	assert RAM(11703) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(11703))))  severity failure;
	assert RAM(11704) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(11704))))  severity failure;
	assert RAM(11705) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(11705))))  severity failure;
	assert RAM(11706) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(11706))))  severity failure;
	assert RAM(11707) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(11707))))  severity failure;
	assert RAM(11708) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(11708))))  severity failure;
	assert RAM(11709) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(11709))))  severity failure;
	assert RAM(11710) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(11710))))  severity failure;
	assert RAM(11711) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(11711))))  severity failure;
	assert RAM(11712) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(11712))))  severity failure;
	assert RAM(11713) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(11713))))  severity failure;
	assert RAM(11714) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(11714))))  severity failure;
	assert RAM(11715) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(11715))))  severity failure;
	assert RAM(11716) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(11716))))  severity failure;
	assert RAM(11717) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(11717))))  severity failure;
	assert RAM(11718) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(11718))))  severity failure;
	assert RAM(11719) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(11719))))  severity failure;
	assert RAM(11720) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(11720))))  severity failure;
	assert RAM(11721) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(11721))))  severity failure;
	assert RAM(11722) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(11722))))  severity failure;
	assert RAM(11723) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(11723))))  severity failure;
	assert RAM(11724) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(11724))))  severity failure;
	assert RAM(11725) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(11725))))  severity failure;
	assert RAM(11726) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(11726))))  severity failure;
	assert RAM(11727) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(11727))))  severity failure;
	assert RAM(11728) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(11728))))  severity failure;
	assert RAM(11729) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(11729))))  severity failure;
	assert RAM(11730) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(11730))))  severity failure;
	assert RAM(11731) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(11731))))  severity failure;
	assert RAM(11732) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(11732))))  severity failure;
	assert RAM(11733) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(11733))))  severity failure;
	assert RAM(11734) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(11734))))  severity failure;
	assert RAM(11735) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(11735))))  severity failure;
	assert RAM(11736) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(11736))))  severity failure;
	assert RAM(11737) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(11737))))  severity failure;
	assert RAM(11738) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(11738))))  severity failure;
	assert RAM(11739) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(11739))))  severity failure;
	assert RAM(11740) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(11740))))  severity failure;
	assert RAM(11741) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(11741))))  severity failure;
	assert RAM(11742) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(11742))))  severity failure;
	assert RAM(11743) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(11743))))  severity failure;
	assert RAM(11744) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(11744))))  severity failure;
	assert RAM(11745) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(11745))))  severity failure;
	assert RAM(11746) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(11746))))  severity failure;
	assert RAM(11747) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(11747))))  severity failure;
	assert RAM(11748) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(11748))))  severity failure;
	assert RAM(11749) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(11749))))  severity failure;
	assert RAM(11750) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(11750))))  severity failure;
	assert RAM(11751) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(11751))))  severity failure;
	assert RAM(11752) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(11752))))  severity failure;
	assert RAM(11753) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(11753))))  severity failure;
	assert RAM(11754) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(11754))))  severity failure;
	assert RAM(11755) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(11755))))  severity failure;
	assert RAM(11756) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(11756))))  severity failure;
	assert RAM(11757) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(11757))))  severity failure;
	assert RAM(11758) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(11758))))  severity failure;
	assert RAM(11759) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(11759))))  severity failure;
	assert RAM(11760) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(11760))))  severity failure;
	assert RAM(11761) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(11761))))  severity failure;
	assert RAM(11762) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(11762))))  severity failure;
	assert RAM(11763) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(11763))))  severity failure;
	assert RAM(11764) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(11764))))  severity failure;
	assert RAM(11765) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(11765))))  severity failure;
	assert RAM(11766) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(11766))))  severity failure;
	assert RAM(11767) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(11767))))  severity failure;
	assert RAM(11768) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(11768))))  severity failure;
	assert RAM(11769) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(11769))))  severity failure;
	assert RAM(11770) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(11770))))  severity failure;
	assert RAM(11771) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(11771))))  severity failure;
	assert RAM(11772) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(11772))))  severity failure;
	assert RAM(11773) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(11773))))  severity failure;
	assert RAM(11774) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(11774))))  severity failure;
	assert RAM(11775) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(11775))))  severity failure;
	assert RAM(11776) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(11776))))  severity failure;
	assert RAM(11777) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(11777))))  severity failure;
	assert RAM(11778) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(11778))))  severity failure;
	assert RAM(11779) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(11779))))  severity failure;
	assert RAM(11780) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(11780))))  severity failure;
	assert RAM(11781) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(11781))))  severity failure;
	assert RAM(11782) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(11782))))  severity failure;
	assert RAM(11783) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(11783))))  severity failure;
	assert RAM(11784) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(11784))))  severity failure;
	assert RAM(11785) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(11785))))  severity failure;
	assert RAM(11786) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(11786))))  severity failure;
	assert RAM(11787) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(11787))))  severity failure;
	assert RAM(11788) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(11788))))  severity failure;
	assert RAM(11789) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(11789))))  severity failure;
	assert RAM(11790) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(11790))))  severity failure;
	assert RAM(11791) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(11791))))  severity failure;
	assert RAM(11792) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(11792))))  severity failure;
	assert RAM(11793) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(11793))))  severity failure;
	assert RAM(11794) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(11794))))  severity failure;
	assert RAM(11795) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(11795))))  severity failure;
	assert RAM(11796) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(11796))))  severity failure;
	assert RAM(11797) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(11797))))  severity failure;
	assert RAM(11798) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(11798))))  severity failure;
	assert RAM(11799) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(11799))))  severity failure;
	assert RAM(11800) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(11800))))  severity failure;
	assert RAM(11801) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(11801))))  severity failure;
	assert RAM(11802) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(11802))))  severity failure;
	assert RAM(11803) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(11803))))  severity failure;
	assert RAM(11804) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(11804))))  severity failure;
	assert RAM(11805) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(11805))))  severity failure;
	assert RAM(11806) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(11806))))  severity failure;
	assert RAM(11807) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(11807))))  severity failure;
	assert RAM(11808) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(11808))))  severity failure;
	assert RAM(11809) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(11809))))  severity failure;
	assert RAM(11810) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(11810))))  severity failure;
	assert RAM(11811) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(11811))))  severity failure;
	assert RAM(11812) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(11812))))  severity failure;
	assert RAM(11813) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(11813))))  severity failure;
	assert RAM(11814) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(11814))))  severity failure;
	assert RAM(11815) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(11815))))  severity failure;
	assert RAM(11816) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(11816))))  severity failure;
	assert RAM(11817) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(11817))))  severity failure;
	assert RAM(11818) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(11818))))  severity failure;
	assert RAM(11819) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(11819))))  severity failure;
	assert RAM(11820) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(11820))))  severity failure;
	assert RAM(11821) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(11821))))  severity failure;
	assert RAM(11822) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(11822))))  severity failure;
	assert RAM(11823) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(11823))))  severity failure;
	assert RAM(11824) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(11824))))  severity failure;
	assert RAM(11825) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(11825))))  severity failure;
	assert RAM(11826) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(11826))))  severity failure;
	assert RAM(11827) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(11827))))  severity failure;
	assert RAM(11828) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(11828))))  severity failure;
	assert RAM(11829) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(11829))))  severity failure;
	assert RAM(11830) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(11830))))  severity failure;
	assert RAM(11831) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(11831))))  severity failure;
	assert RAM(11832) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(11832))))  severity failure;
	assert RAM(11833) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(11833))))  severity failure;
	assert RAM(11834) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(11834))))  severity failure;
	assert RAM(11835) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(11835))))  severity failure;
	assert RAM(11836) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(11836))))  severity failure;
	assert RAM(11837) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(11837))))  severity failure;
	assert RAM(11838) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(11838))))  severity failure;
	assert RAM(11839) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(11839))))  severity failure;
	assert RAM(11840) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(11840))))  severity failure;
	assert RAM(11841) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(11841))))  severity failure;
	assert RAM(11842) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(11842))))  severity failure;
	assert RAM(11843) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(11843))))  severity failure;
	assert RAM(11844) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(11844))))  severity failure;
	assert RAM(11845) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(11845))))  severity failure;
	assert RAM(11846) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(11846))))  severity failure;
	assert RAM(11847) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(11847))))  severity failure;
	assert RAM(11848) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(11848))))  severity failure;
	assert RAM(11849) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(11849))))  severity failure;
	assert RAM(11850) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(11850))))  severity failure;
	assert RAM(11851) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(11851))))  severity failure;
	assert RAM(11852) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(11852))))  severity failure;
	assert RAM(11853) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(11853))))  severity failure;
	assert RAM(11854) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(11854))))  severity failure;
	assert RAM(11855) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(11855))))  severity failure;
	assert RAM(11856) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(11856))))  severity failure;
	assert RAM(11857) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(11857))))  severity failure;
	assert RAM(11858) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(11858))))  severity failure;
	assert RAM(11859) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(11859))))  severity failure;
	assert RAM(11860) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(11860))))  severity failure;
	assert RAM(11861) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(11861))))  severity failure;
	assert RAM(11862) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(11862))))  severity failure;
	assert RAM(11863) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(11863))))  severity failure;
	assert RAM(11864) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(11864))))  severity failure;
	assert RAM(11865) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(11865))))  severity failure;
	assert RAM(11866) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(11866))))  severity failure;
	assert RAM(11867) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(11867))))  severity failure;
	assert RAM(11868) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(11868))))  severity failure;
	assert RAM(11869) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(11869))))  severity failure;
	assert RAM(11870) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(11870))))  severity failure;
	assert RAM(11871) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(11871))))  severity failure;
	assert RAM(11872) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(11872))))  severity failure;
	assert RAM(11873) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(11873))))  severity failure;
	assert RAM(11874) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(11874))))  severity failure;
	assert RAM(11875) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(11875))))  severity failure;
	assert RAM(11876) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(11876))))  severity failure;
	assert RAM(11877) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(11877))))  severity failure;
	assert RAM(11878) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(11878))))  severity failure;
	assert RAM(11879) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(11879))))  severity failure;
	assert RAM(11880) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(11880))))  severity failure;
	assert RAM(11881) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(11881))))  severity failure;
	assert RAM(11882) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(11882))))  severity failure;
	assert RAM(11883) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(11883))))  severity failure;
	assert RAM(11884) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(11884))))  severity failure;
	assert RAM(11885) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(11885))))  severity failure;
	assert RAM(11886) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(11886))))  severity failure;
	assert RAM(11887) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(11887))))  severity failure;
	assert RAM(11888) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(11888))))  severity failure;
	assert RAM(11889) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(11889))))  severity failure;
	assert RAM(11890) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(11890))))  severity failure;
	assert RAM(11891) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(11891))))  severity failure;
	assert RAM(11892) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(11892))))  severity failure;
	assert RAM(11893) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(11893))))  severity failure;
	assert RAM(11894) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(11894))))  severity failure;
	assert RAM(11895) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(11895))))  severity failure;
	assert RAM(11896) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(11896))))  severity failure;
	assert RAM(11897) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(11897))))  severity failure;
	assert RAM(11898) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(11898))))  severity failure;
	assert RAM(11899) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(11899))))  severity failure;
	assert RAM(11900) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(11900))))  severity failure;
	assert RAM(11901) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(11901))))  severity failure;
	assert RAM(11902) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(11902))))  severity failure;
	assert RAM(11903) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(11903))))  severity failure;
	assert RAM(11904) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(11904))))  severity failure;
	assert RAM(11905) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(11905))))  severity failure;
	assert RAM(11906) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(11906))))  severity failure;
	assert RAM(11907) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(11907))))  severity failure;
	assert RAM(11908) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(11908))))  severity failure;
	assert RAM(11909) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(11909))))  severity failure;
	assert RAM(11910) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(11910))))  severity failure;
	assert RAM(11911) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(11911))))  severity failure;
	assert RAM(11912) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(11912))))  severity failure;
	assert RAM(11913) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(11913))))  severity failure;
	assert RAM(11914) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(11914))))  severity failure;
	assert RAM(11915) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(11915))))  severity failure;
	assert RAM(11916) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(11916))))  severity failure;
	assert RAM(11917) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(11917))))  severity failure;
	assert RAM(11918) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(11918))))  severity failure;
	assert RAM(11919) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(11919))))  severity failure;
	assert RAM(11920) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(11920))))  severity failure;
	assert RAM(11921) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(11921))))  severity failure;
	assert RAM(11922) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(11922))))  severity failure;
	assert RAM(11923) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(11923))))  severity failure;
	assert RAM(11924) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(11924))))  severity failure;
	assert RAM(11925) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(11925))))  severity failure;
	assert RAM(11926) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(11926))))  severity failure;
	assert RAM(11927) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(11927))))  severity failure;
	assert RAM(11928) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(11928))))  severity failure;
	assert RAM(11929) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(11929))))  severity failure;
	assert RAM(11930) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(11930))))  severity failure;
	assert RAM(11931) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(11931))))  severity failure;
	assert RAM(11932) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(11932))))  severity failure;
	assert RAM(11933) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(11933))))  severity failure;
	assert RAM(11934) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(11934))))  severity failure;
	assert RAM(11935) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(11935))))  severity failure;
	assert RAM(11936) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(11936))))  severity failure;
	assert RAM(11937) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(11937))))  severity failure;
	assert RAM(11938) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(11938))))  severity failure;
	assert RAM(11939) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(11939))))  severity failure;
	assert RAM(11940) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(11940))))  severity failure;
	assert RAM(11941) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(11941))))  severity failure;
	assert RAM(11942) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(11942))))  severity failure;
	assert RAM(11943) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(11943))))  severity failure;
	assert RAM(11944) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(11944))))  severity failure;
	assert RAM(11945) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(11945))))  severity failure;
	assert RAM(11946) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(11946))))  severity failure;
	assert RAM(11947) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(11947))))  severity failure;
	assert RAM(11948) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(11948))))  severity failure;
	assert RAM(11949) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(11949))))  severity failure;
	assert RAM(11950) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(11950))))  severity failure;
	assert RAM(11951) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(11951))))  severity failure;
	assert RAM(11952) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(11952))))  severity failure;
	assert RAM(11953) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(11953))))  severity failure;
	assert RAM(11954) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(11954))))  severity failure;
	assert RAM(11955) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(11955))))  severity failure;
	assert RAM(11956) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(11956))))  severity failure;
	assert RAM(11957) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(11957))))  severity failure;
	assert RAM(11958) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(11958))))  severity failure;
	assert RAM(11959) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(11959))))  severity failure;
	assert RAM(11960) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(11960))))  severity failure;
	assert RAM(11961) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(11961))))  severity failure;
	assert RAM(11962) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(11962))))  severity failure;
	assert RAM(11963) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(11963))))  severity failure;
	assert RAM(11964) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(11964))))  severity failure;
	assert RAM(11965) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(11965))))  severity failure;
	assert RAM(11966) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(11966))))  severity failure;
	assert RAM(11967) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(11967))))  severity failure;
	assert RAM(11968) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(11968))))  severity failure;
	assert RAM(11969) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(11969))))  severity failure;
	assert RAM(11970) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(11970))))  severity failure;
	assert RAM(11971) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(11971))))  severity failure;
	assert RAM(11972) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(11972))))  severity failure;
	assert RAM(11973) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(11973))))  severity failure;
	assert RAM(11974) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(11974))))  severity failure;
	assert RAM(11975) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(11975))))  severity failure;
	assert RAM(11976) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(11976))))  severity failure;
	assert RAM(11977) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(11977))))  severity failure;
	assert RAM(11978) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(11978))))  severity failure;
	assert RAM(11979) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(11979))))  severity failure;
	assert RAM(11980) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(11980))))  severity failure;
	assert RAM(11981) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(11981))))  severity failure;
	assert RAM(11982) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(11982))))  severity failure;
	assert RAM(11983) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(11983))))  severity failure;
	assert RAM(11984) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(11984))))  severity failure;
	assert RAM(11985) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(11985))))  severity failure;
	assert RAM(11986) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(11986))))  severity failure;
	assert RAM(11987) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(11987))))  severity failure;
	assert RAM(11988) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(11988))))  severity failure;
	assert RAM(11989) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(11989))))  severity failure;
	assert RAM(11990) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(11990))))  severity failure;
	assert RAM(11991) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(11991))))  severity failure;
	assert RAM(11992) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(11992))))  severity failure;
	assert RAM(11993) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(11993))))  severity failure;
	assert RAM(11994) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(11994))))  severity failure;
	assert RAM(11995) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(11995))))  severity failure;
	assert RAM(11996) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(11996))))  severity failure;
	assert RAM(11997) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(11997))))  severity failure;
	assert RAM(11998) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(11998))))  severity failure;
	assert RAM(11999) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(11999))))  severity failure;
	assert RAM(12000) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(12000))))  severity failure;
	assert RAM(12001) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(12001))))  severity failure;
	assert RAM(12002) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(12002))))  severity failure;
	assert RAM(12003) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(12003))))  severity failure;
	assert RAM(12004) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(12004))))  severity failure;
	assert RAM(12005) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(12005))))  severity failure;
	assert RAM(12006) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(12006))))  severity failure;
	assert RAM(12007) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(12007))))  severity failure;
	assert RAM(12008) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(12008))))  severity failure;
	assert RAM(12009) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(12009))))  severity failure;
	assert RAM(12010) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(12010))))  severity failure;
	assert RAM(12011) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(12011))))  severity failure;
	assert RAM(12012) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(12012))))  severity failure;
	assert RAM(12013) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(12013))))  severity failure;
	assert RAM(12014) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(12014))))  severity failure;
	assert RAM(12015) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(12015))))  severity failure;
	assert RAM(12016) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(12016))))  severity failure;
	assert RAM(12017) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(12017))))  severity failure;
	assert RAM(12018) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(12018))))  severity failure;
	assert RAM(12019) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(12019))))  severity failure;
	assert RAM(12020) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(12020))))  severity failure;
	assert RAM(12021) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(12021))))  severity failure;
	assert RAM(12022) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(12022))))  severity failure;
	assert RAM(12023) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(12023))))  severity failure;
	assert RAM(12024) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(12024))))  severity failure;
	assert RAM(12025) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(12025))))  severity failure;
	assert RAM(12026) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(12026))))  severity failure;
	assert RAM(12027) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(12027))))  severity failure;
	assert RAM(12028) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(12028))))  severity failure;
	assert RAM(12029) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(12029))))  severity failure;
	assert RAM(12030) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(12030))))  severity failure;
	assert RAM(12031) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(12031))))  severity failure;
	assert RAM(12032) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(12032))))  severity failure;
	assert RAM(12033) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(12033))))  severity failure;
	assert RAM(12034) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(12034))))  severity failure;
	assert RAM(12035) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(12035))))  severity failure;
	assert RAM(12036) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(12036))))  severity failure;
	assert RAM(12037) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(12037))))  severity failure;
	assert RAM(12038) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(12038))))  severity failure;
	assert RAM(12039) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(12039))))  severity failure;
	assert RAM(12040) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(12040))))  severity failure;
	assert RAM(12041) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(12041))))  severity failure;
	assert RAM(12042) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(12042))))  severity failure;
	assert RAM(12043) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(12043))))  severity failure;
	assert RAM(12044) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(12044))))  severity failure;
	assert RAM(12045) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(12045))))  severity failure;
	assert RAM(12046) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(12046))))  severity failure;
	assert RAM(12047) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(12047))))  severity failure;
	assert RAM(12048) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(12048))))  severity failure;
	assert RAM(12049) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(12049))))  severity failure;
	assert RAM(12050) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(12050))))  severity failure;
	assert RAM(12051) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(12051))))  severity failure;
	assert RAM(12052) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(12052))))  severity failure;
	assert RAM(12053) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(12053))))  severity failure;
	assert RAM(12054) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(12054))))  severity failure;
	assert RAM(12055) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(12055))))  severity failure;
	assert RAM(12056) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(12056))))  severity failure;
	assert RAM(12057) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(12057))))  severity failure;
	assert RAM(12058) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(12058))))  severity failure;
	assert RAM(12059) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(12059))))  severity failure;
	assert RAM(12060) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(12060))))  severity failure;
	assert RAM(12061) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(12061))))  severity failure;
	assert RAM(12062) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(12062))))  severity failure;
	assert RAM(12063) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(12063))))  severity failure;
	assert RAM(12064) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(12064))))  severity failure;
	assert RAM(12065) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(12065))))  severity failure;
	assert RAM(12066) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(12066))))  severity failure;
	assert RAM(12067) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(12067))))  severity failure;
	assert RAM(12068) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(12068))))  severity failure;
	assert RAM(12069) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(12069))))  severity failure;
	assert RAM(12070) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(12070))))  severity failure;
	assert RAM(12071) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(12071))))  severity failure;
	assert RAM(12072) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(12072))))  severity failure;
	assert RAM(12073) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(12073))))  severity failure;
	assert RAM(12074) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(12074))))  severity failure;
	assert RAM(12075) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(12075))))  severity failure;
	assert RAM(12076) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(12076))))  severity failure;
	assert RAM(12077) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(12077))))  severity failure;
	assert RAM(12078) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(12078))))  severity failure;
	assert RAM(12079) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(12079))))  severity failure;
	assert RAM(12080) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(12080))))  severity failure;
	assert RAM(12081) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(12081))))  severity failure;
	assert RAM(12082) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(12082))))  severity failure;
	assert RAM(12083) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(12083))))  severity failure;
	assert RAM(12084) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(12084))))  severity failure;
	assert RAM(12085) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(12085))))  severity failure;
	assert RAM(12086) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(12086))))  severity failure;
	assert RAM(12087) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(12087))))  severity failure;
	assert RAM(12088) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(12088))))  severity failure;
	assert RAM(12089) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(12089))))  severity failure;
	assert RAM(12090) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(12090))))  severity failure;
	assert RAM(12091) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(12091))))  severity failure;
	assert RAM(12092) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(12092))))  severity failure;
	assert RAM(12093) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(12093))))  severity failure;
	assert RAM(12094) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(12094))))  severity failure;
	assert RAM(12095) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(12095))))  severity failure;
	assert RAM(12096) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(12096))))  severity failure;
	assert RAM(12097) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(12097))))  severity failure;
	assert RAM(12098) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(12098))))  severity failure;
	assert RAM(12099) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(12099))))  severity failure;
	assert RAM(12100) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(12100))))  severity failure;
	assert RAM(12101) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(12101))))  severity failure;
	assert RAM(12102) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(12102))))  severity failure;
	assert RAM(12103) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(12103))))  severity failure;
	assert RAM(12104) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(12104))))  severity failure;
	assert RAM(12105) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(12105))))  severity failure;
	assert RAM(12106) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(12106))))  severity failure;
	assert RAM(12107) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(12107))))  severity failure;
	assert RAM(12108) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(12108))))  severity failure;
	assert RAM(12109) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(12109))))  severity failure;
	assert RAM(12110) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(12110))))  severity failure;
	assert RAM(12111) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(12111))))  severity failure;
	assert RAM(12112) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(12112))))  severity failure;
	assert RAM(12113) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(12113))))  severity failure;
	assert RAM(12114) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(12114))))  severity failure;
	assert RAM(12115) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(12115))))  severity failure;
	assert RAM(12116) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(12116))))  severity failure;
	assert RAM(12117) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(12117))))  severity failure;
	assert RAM(12118) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(12118))))  severity failure;
	assert RAM(12119) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(12119))))  severity failure;
	assert RAM(12120) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(12120))))  severity failure;
	assert RAM(12121) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(12121))))  severity failure;
	assert RAM(12122) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(12122))))  severity failure;
	assert RAM(12123) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(12123))))  severity failure;
	assert RAM(12124) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(12124))))  severity failure;
	assert RAM(12125) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(12125))))  severity failure;
	assert RAM(12126) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(12126))))  severity failure;
	assert RAM(12127) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(12127))))  severity failure;
	assert RAM(12128) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(12128))))  severity failure;
	assert RAM(12129) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(12129))))  severity failure;
	assert RAM(12130) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(12130))))  severity failure;
	assert RAM(12131) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(12131))))  severity failure;
	assert RAM(12132) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(12132))))  severity failure;
	assert RAM(12133) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(12133))))  severity failure;
	assert RAM(12134) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(12134))))  severity failure;
	assert RAM(12135) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(12135))))  severity failure;
	assert RAM(12136) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(12136))))  severity failure;
	assert RAM(12137) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(12137))))  severity failure;
	assert RAM(12138) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(12138))))  severity failure;
	assert RAM(12139) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(12139))))  severity failure;
	assert RAM(12140) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(12140))))  severity failure;
	assert RAM(12141) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(12141))))  severity failure;
	assert RAM(12142) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(12142))))  severity failure;
	assert RAM(12143) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(12143))))  severity failure;
	assert RAM(12144) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(12144))))  severity failure;
	assert RAM(12145) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(12145))))  severity failure;
	assert RAM(12146) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(12146))))  severity failure;
	assert RAM(12147) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(12147))))  severity failure;
	assert RAM(12148) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(12148))))  severity failure;
	assert RAM(12149) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(12149))))  severity failure;
	assert RAM(12150) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(12150))))  severity failure;
	assert RAM(12151) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(12151))))  severity failure;
	assert RAM(12152) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(12152))))  severity failure;
	assert RAM(12153) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(12153))))  severity failure;
	assert RAM(12154) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(12154))))  severity failure;
	assert RAM(12155) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(12155))))  severity failure;
	assert RAM(12156) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(12156))))  severity failure;
	assert RAM(12157) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(12157))))  severity failure;
	assert RAM(12158) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(12158))))  severity failure;
	assert RAM(12159) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(12159))))  severity failure;
	assert RAM(12160) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(12160))))  severity failure;
	assert RAM(12161) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(12161))))  severity failure;
	assert RAM(12162) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(12162))))  severity failure;
	assert RAM(12163) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(12163))))  severity failure;
	assert RAM(12164) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(12164))))  severity failure;
	assert RAM(12165) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(12165))))  severity failure;
	assert RAM(12166) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(12166))))  severity failure;
	assert RAM(12167) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(12167))))  severity failure;
	assert RAM(12168) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(12168))))  severity failure;
	assert RAM(12169) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(12169))))  severity failure;
	assert RAM(12170) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(12170))))  severity failure;
	assert RAM(12171) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(12171))))  severity failure;
	assert RAM(12172) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(12172))))  severity failure;
	assert RAM(12173) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(12173))))  severity failure;
	assert RAM(12174) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(12174))))  severity failure;
	assert RAM(12175) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(12175))))  severity failure;
	assert RAM(12176) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(12176))))  severity failure;
	assert RAM(12177) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(12177))))  severity failure;
	assert RAM(12178) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(12178))))  severity failure;
	assert RAM(12179) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(12179))))  severity failure;
	assert RAM(12180) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(12180))))  severity failure;
	assert RAM(12181) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(12181))))  severity failure;
	assert RAM(12182) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(12182))))  severity failure;
	assert RAM(12183) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(12183))))  severity failure;
	assert RAM(12184) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(12184))))  severity failure;
	assert RAM(12185) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(12185))))  severity failure;
	assert RAM(12186) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(12186))))  severity failure;
	assert RAM(12187) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(12187))))  severity failure;
	assert RAM(12188) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(12188))))  severity failure;
	assert RAM(12189) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(12189))))  severity failure;
	assert RAM(12190) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(12190))))  severity failure;
	assert RAM(12191) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(12191))))  severity failure;
	assert RAM(12192) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(12192))))  severity failure;
	assert RAM(12193) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(12193))))  severity failure;
	assert RAM(12194) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(12194))))  severity failure;
	assert RAM(12195) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(12195))))  severity failure;
	assert RAM(12196) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(12196))))  severity failure;
	assert RAM(12197) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(12197))))  severity failure;
	assert RAM(12198) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(12198))))  severity failure;
	assert RAM(12199) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(12199))))  severity failure;
	assert RAM(12200) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(12200))))  severity failure;
	assert RAM(12201) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(12201))))  severity failure;
	assert RAM(12202) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(12202))))  severity failure;
	assert RAM(12203) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(12203))))  severity failure;
	assert RAM(12204) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(12204))))  severity failure;
	assert RAM(12205) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(12205))))  severity failure;
	assert RAM(12206) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(12206))))  severity failure;
	assert RAM(12207) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(12207))))  severity failure;
	assert RAM(12208) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(12208))))  severity failure;
	assert RAM(12209) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(12209))))  severity failure;
	assert RAM(12210) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(12210))))  severity failure;
	assert RAM(12211) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(12211))))  severity failure;
	assert RAM(12212) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(12212))))  severity failure;
	assert RAM(12213) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(12213))))  severity failure;
	assert RAM(12214) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(12214))))  severity failure;
	assert RAM(12215) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(12215))))  severity failure;
	assert RAM(12216) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(12216))))  severity failure;
	assert RAM(12217) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(12217))))  severity failure;
	assert RAM(12218) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(12218))))  severity failure;
	assert RAM(12219) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(12219))))  severity failure;
	assert RAM(12220) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(12220))))  severity failure;
	assert RAM(12221) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(12221))))  severity failure;
	assert RAM(12222) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(12222))))  severity failure;
	assert RAM(12223) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(12223))))  severity failure;
	assert RAM(12224) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(12224))))  severity failure;
	assert RAM(12225) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(12225))))  severity failure;
	assert RAM(12226) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(12226))))  severity failure;
	assert RAM(12227) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(12227))))  severity failure;
	assert RAM(12228) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(12228))))  severity failure;
	assert RAM(12229) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(12229))))  severity failure;
	assert RAM(12230) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(12230))))  severity failure;
	assert RAM(12231) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(12231))))  severity failure;
	assert RAM(12232) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(12232))))  severity failure;
	assert RAM(12233) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(12233))))  severity failure;
	assert RAM(12234) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(12234))))  severity failure;
	assert RAM(12235) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(12235))))  severity failure;
	assert RAM(12236) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(12236))))  severity failure;
	assert RAM(12237) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(12237))))  severity failure;
	assert RAM(12238) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(12238))))  severity failure;
	assert RAM(12239) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(12239))))  severity failure;
	assert RAM(12240) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(12240))))  severity failure;
	assert RAM(12241) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(12241))))  severity failure;
	assert RAM(12242) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(12242))))  severity failure;
	assert RAM(12243) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(12243))))  severity failure;
	assert RAM(12244) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(12244))))  severity failure;
	assert RAM(12245) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(12245))))  severity failure;
	assert RAM(12246) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(12246))))  severity failure;
	assert RAM(12247) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(12247))))  severity failure;
	assert RAM(12248) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(12248))))  severity failure;
	assert RAM(12249) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(12249))))  severity failure;
	assert RAM(12250) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(12250))))  severity failure;
	assert RAM(12251) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(12251))))  severity failure;
	assert RAM(12252) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(12252))))  severity failure;
	assert RAM(12253) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(12253))))  severity failure;
	assert RAM(12254) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(12254))))  severity failure;
	assert RAM(12255) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(12255))))  severity failure;
	assert RAM(12256) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(12256))))  severity failure;
	assert RAM(12257) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(12257))))  severity failure;
	assert RAM(12258) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(12258))))  severity failure;
	assert RAM(12259) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(12259))))  severity failure;
	assert RAM(12260) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(12260))))  severity failure;
	assert RAM(12261) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(12261))))  severity failure;
	assert RAM(12262) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(12262))))  severity failure;
	assert RAM(12263) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(12263))))  severity failure;
	assert RAM(12264) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(12264))))  severity failure;
	assert RAM(12265) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(12265))))  severity failure;
	assert RAM(12266) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(12266))))  severity failure;
	assert RAM(12267) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(12267))))  severity failure;
	assert RAM(12268) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(12268))))  severity failure;
	assert RAM(12269) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(12269))))  severity failure;
	assert RAM(12270) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(12270))))  severity failure;
	assert RAM(12271) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(12271))))  severity failure;
	assert RAM(12272) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(12272))))  severity failure;
	assert RAM(12273) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(12273))))  severity failure;
	assert RAM(12274) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(12274))))  severity failure;
	assert RAM(12275) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(12275))))  severity failure;
	assert RAM(12276) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(12276))))  severity failure;
	assert RAM(12277) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(12277))))  severity failure;
	assert RAM(12278) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(12278))))  severity failure;
	assert RAM(12279) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(12279))))  severity failure;
	assert RAM(12280) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(12280))))  severity failure;
	assert RAM(12281) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(12281))))  severity failure;
	assert RAM(12282) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(12282))))  severity failure;
	assert RAM(12283) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(12283))))  severity failure;
	assert RAM(12284) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(12284))))  severity failure;
	assert RAM(12285) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(12285))))  severity failure;
	assert RAM(12286) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(12286))))  severity failure;
	assert RAM(12287) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(12287))))  severity failure;
	assert RAM(12288) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(12288))))  severity failure;
	assert RAM(12289) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(12289))))  severity failure;
	assert RAM(12290) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(12290))))  severity failure;
	assert RAM(12291) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(12291))))  severity failure;
	assert RAM(12292) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(12292))))  severity failure;
	assert RAM(12293) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(12293))))  severity failure;
	assert RAM(12294) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(12294))))  severity failure;
	assert RAM(12295) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(12295))))  severity failure;
	assert RAM(12296) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(12296))))  severity failure;
	assert RAM(12297) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(12297))))  severity failure;
	assert RAM(12298) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(12298))))  severity failure;
	assert RAM(12299) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(12299))))  severity failure;
	assert RAM(12300) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(12300))))  severity failure;
	assert RAM(12301) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(12301))))  severity failure;
	assert RAM(12302) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(12302))))  severity failure;
	assert RAM(12303) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(12303))))  severity failure;
	assert RAM(12304) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(12304))))  severity failure;
	assert RAM(12305) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(12305))))  severity failure;
	assert RAM(12306) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(12306))))  severity failure;
	assert RAM(12307) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(12307))))  severity failure;
	assert RAM(12308) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(12308))))  severity failure;
	assert RAM(12309) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(12309))))  severity failure;
	assert RAM(12310) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(12310))))  severity failure;
	assert RAM(12311) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(12311))))  severity failure;
	assert RAM(12312) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(12312))))  severity failure;
	assert RAM(12313) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(12313))))  severity failure;
	assert RAM(12314) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(12314))))  severity failure;
	assert RAM(12315) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(12315))))  severity failure;
	assert RAM(12316) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(12316))))  severity failure;
	assert RAM(12317) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(12317))))  severity failure;
	assert RAM(12318) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(12318))))  severity failure;
	assert RAM(12319) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(12319))))  severity failure;
	assert RAM(12320) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(12320))))  severity failure;
	assert RAM(12321) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(12321))))  severity failure;
	assert RAM(12322) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(12322))))  severity failure;
	assert RAM(12323) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(12323))))  severity failure;
	assert RAM(12324) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(12324))))  severity failure;
	assert RAM(12325) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(12325))))  severity failure;
	assert RAM(12326) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(12326))))  severity failure;
	assert RAM(12327) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(12327))))  severity failure;
	assert RAM(12328) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(12328))))  severity failure;
	assert RAM(12329) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(12329))))  severity failure;
	assert RAM(12330) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(12330))))  severity failure;
	assert RAM(12331) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(12331))))  severity failure;
	assert RAM(12332) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(12332))))  severity failure;
	assert RAM(12333) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(12333))))  severity failure;
	assert RAM(12334) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(12334))))  severity failure;
	assert RAM(12335) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(12335))))  severity failure;
	assert RAM(12336) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(12336))))  severity failure;
	assert RAM(12337) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(12337))))  severity failure;
	assert RAM(12338) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(12338))))  severity failure;
	assert RAM(12339) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(12339))))  severity failure;
	assert RAM(12340) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(12340))))  severity failure;
	assert RAM(12341) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(12341))))  severity failure;
	assert RAM(12342) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(12342))))  severity failure;
	assert RAM(12343) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(12343))))  severity failure;
	assert RAM(12344) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(12344))))  severity failure;
	assert RAM(12345) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(12345))))  severity failure;
	assert RAM(12346) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(12346))))  severity failure;
	assert RAM(12347) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(12347))))  severity failure;
	assert RAM(12348) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(12348))))  severity failure;
	assert RAM(12349) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(12349))))  severity failure;
	assert RAM(12350) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(12350))))  severity failure;
	assert RAM(12351) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(12351))))  severity failure;
	assert RAM(12352) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(12352))))  severity failure;
	assert RAM(12353) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(12353))))  severity failure;
	assert RAM(12354) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(12354))))  severity failure;
	assert RAM(12355) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(12355))))  severity failure;
	assert RAM(12356) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(12356))))  severity failure;
	assert RAM(12357) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(12357))))  severity failure;
	assert RAM(12358) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(12358))))  severity failure;
	assert RAM(12359) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(12359))))  severity failure;
	assert RAM(12360) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(12360))))  severity failure;
	assert RAM(12361) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(12361))))  severity failure;
	assert RAM(12362) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(12362))))  severity failure;
	assert RAM(12363) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(12363))))  severity failure;
	assert RAM(12364) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(12364))))  severity failure;
	assert RAM(12365) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(12365))))  severity failure;
	assert RAM(12366) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(12366))))  severity failure;
	assert RAM(12367) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(12367))))  severity failure;
	assert RAM(12368) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(12368))))  severity failure;
	assert RAM(12369) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(12369))))  severity failure;
	assert RAM(12370) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(12370))))  severity failure;
	assert RAM(12371) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(12371))))  severity failure;
	assert RAM(12372) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(12372))))  severity failure;
	assert RAM(12373) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(12373))))  severity failure;
	assert RAM(12374) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(12374))))  severity failure;
	assert RAM(12375) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(12375))))  severity failure;
	assert RAM(12376) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(12376))))  severity failure;
	assert RAM(12377) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(12377))))  severity failure;
	assert RAM(12378) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(12378))))  severity failure;
	assert RAM(12379) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(12379))))  severity failure;
	assert RAM(12380) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(12380))))  severity failure;
	assert RAM(12381) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(12381))))  severity failure;
	assert RAM(12382) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(12382))))  severity failure;
	assert RAM(12383) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(12383))))  severity failure;
	assert RAM(12384) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(12384))))  severity failure;
	assert RAM(12385) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(12385))))  severity failure;
	assert RAM(12386) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(12386))))  severity failure;
	assert RAM(12387) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(12387))))  severity failure;
	assert RAM(12388) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(12388))))  severity failure;
	assert RAM(12389) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(12389))))  severity failure;
	assert RAM(12390) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(12390))))  severity failure;
	assert RAM(12391) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(12391))))  severity failure;
	assert RAM(12392) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(12392))))  severity failure;
	assert RAM(12393) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(12393))))  severity failure;
	assert RAM(12394) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(12394))))  severity failure;
	assert RAM(12395) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(12395))))  severity failure;
	assert RAM(12396) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(12396))))  severity failure;
	assert RAM(12397) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(12397))))  severity failure;
	assert RAM(12398) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(12398))))  severity failure;
	assert RAM(12399) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(12399))))  severity failure;
	assert RAM(12400) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(12400))))  severity failure;
	assert RAM(12401) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(12401))))  severity failure;
	assert RAM(12402) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(12402))))  severity failure;
	assert RAM(12403) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(12403))))  severity failure;
	assert RAM(12404) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(12404))))  severity failure;
	assert RAM(12405) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(12405))))  severity failure;
	assert RAM(12406) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(12406))))  severity failure;
	assert RAM(12407) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(12407))))  severity failure;
	assert RAM(12408) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(12408))))  severity failure;
	assert RAM(12409) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(12409))))  severity failure;
	assert RAM(12410) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(12410))))  severity failure;
	assert RAM(12411) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(12411))))  severity failure;
	assert RAM(12412) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(12412))))  severity failure;
	assert RAM(12413) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(12413))))  severity failure;
	assert RAM(12414) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(12414))))  severity failure;
	assert RAM(12415) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(12415))))  severity failure;
	assert RAM(12416) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(12416))))  severity failure;
	assert RAM(12417) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(12417))))  severity failure;
	assert RAM(12418) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(12418))))  severity failure;
	assert RAM(12419) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(12419))))  severity failure;
	assert RAM(12420) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(12420))))  severity failure;
	assert RAM(12421) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(12421))))  severity failure;
	assert RAM(12422) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(12422))))  severity failure;
	assert RAM(12423) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(12423))))  severity failure;
	assert RAM(12424) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(12424))))  severity failure;
	assert RAM(12425) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(12425))))  severity failure;
	assert RAM(12426) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(12426))))  severity failure;
	assert RAM(12427) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(12427))))  severity failure;
	assert RAM(12428) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(12428))))  severity failure;
	assert RAM(12429) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(12429))))  severity failure;
	assert RAM(12430) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(12430))))  severity failure;
	assert RAM(12431) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(12431))))  severity failure;
	assert RAM(12432) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(12432))))  severity failure;
	assert RAM(12433) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(12433))))  severity failure;
	assert RAM(12434) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(12434))))  severity failure;
	assert RAM(12435) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(12435))))  severity failure;
	assert RAM(12436) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(12436))))  severity failure;
	assert RAM(12437) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(12437))))  severity failure;
	assert RAM(12438) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(12438))))  severity failure;
	assert RAM(12439) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(12439))))  severity failure;
	assert RAM(12440) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(12440))))  severity failure;
	assert RAM(12441) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(12441))))  severity failure;
	assert RAM(12442) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(12442))))  severity failure;
	assert RAM(12443) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(12443))))  severity failure;
	assert RAM(12444) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(12444))))  severity failure;
	assert RAM(12445) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(12445))))  severity failure;
	assert RAM(12446) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(12446))))  severity failure;
	assert RAM(12447) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(12447))))  severity failure;
	assert RAM(12448) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(12448))))  severity failure;
	assert RAM(12449) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(12449))))  severity failure;
	assert RAM(12450) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(12450))))  severity failure;
	assert RAM(12451) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(12451))))  severity failure;
	assert RAM(12452) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(12452))))  severity failure;
	assert RAM(12453) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(12453))))  severity failure;
	assert RAM(12454) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(12454))))  severity failure;
	assert RAM(12455) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(12455))))  severity failure;
	assert RAM(12456) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(12456))))  severity failure;
	assert RAM(12457) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(12457))))  severity failure;
	assert RAM(12458) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(12458))))  severity failure;
	assert RAM(12459) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(12459))))  severity failure;
	assert RAM(12460) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(12460))))  severity failure;
	assert RAM(12461) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(12461))))  severity failure;
	assert RAM(12462) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(12462))))  severity failure;
	assert RAM(12463) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(12463))))  severity failure;
	assert RAM(12464) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(12464))))  severity failure;
	assert RAM(12465) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(12465))))  severity failure;
	assert RAM(12466) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(12466))))  severity failure;
	assert RAM(12467) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(12467))))  severity failure;
	assert RAM(12468) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(12468))))  severity failure;
	assert RAM(12469) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(12469))))  severity failure;
	assert RAM(12470) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(12470))))  severity failure;
	assert RAM(12471) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(12471))))  severity failure;
	assert RAM(12472) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(12472))))  severity failure;
	assert RAM(12473) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(12473))))  severity failure;
	assert RAM(12474) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(12474))))  severity failure;
	assert RAM(12475) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(12475))))  severity failure;
	assert RAM(12476) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(12476))))  severity failure;
	assert RAM(12477) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(12477))))  severity failure;
	assert RAM(12478) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(12478))))  severity failure;
	assert RAM(12479) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(12479))))  severity failure;
	assert RAM(12480) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(12480))))  severity failure;
	assert RAM(12481) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(12481))))  severity failure;
	assert RAM(12482) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(12482))))  severity failure;
	assert RAM(12483) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(12483))))  severity failure;
	assert RAM(12484) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(12484))))  severity failure;
	assert RAM(12485) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(12485))))  severity failure;
	assert RAM(12486) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(12486))))  severity failure;
	assert RAM(12487) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(12487))))  severity failure;
	assert RAM(12488) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(12488))))  severity failure;
	assert RAM(12489) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(12489))))  severity failure;
	assert RAM(12490) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(12490))))  severity failure;
	assert RAM(12491) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(12491))))  severity failure;
	assert RAM(12492) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(12492))))  severity failure;
	assert RAM(12493) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(12493))))  severity failure;
	assert RAM(12494) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(12494))))  severity failure;
	assert RAM(12495) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(12495))))  severity failure;
	assert RAM(12496) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(12496))))  severity failure;
	assert RAM(12497) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(12497))))  severity failure;
	assert RAM(12498) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(12498))))  severity failure;
	assert RAM(12499) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(12499))))  severity failure;
	assert RAM(12500) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(12500))))  severity failure;
	assert RAM(12501) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(12501))))  severity failure;
	assert RAM(12502) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(12502))))  severity failure;
	assert RAM(12503) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(12503))))  severity failure;
	assert RAM(12504) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(12504))))  severity failure;
	assert RAM(12505) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(12505))))  severity failure;
	assert RAM(12506) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(12506))))  severity failure;
	assert RAM(12507) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(12507))))  severity failure;
	assert RAM(12508) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(12508))))  severity failure;
	assert RAM(12509) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(12509))))  severity failure;
	assert RAM(12510) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(12510))))  severity failure;
	assert RAM(12511) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(12511))))  severity failure;
	assert RAM(12512) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(12512))))  severity failure;
	assert RAM(12513) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(12513))))  severity failure;
	assert RAM(12514) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(12514))))  severity failure;
	assert RAM(12515) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(12515))))  severity failure;
	assert RAM(12516) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(12516))))  severity failure;
	assert RAM(12517) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(12517))))  severity failure;
	assert RAM(12518) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(12518))))  severity failure;
	assert RAM(12519) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(12519))))  severity failure;
	assert RAM(12520) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(12520))))  severity failure;
	assert RAM(12521) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(12521))))  severity failure;
	assert RAM(12522) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(12522))))  severity failure;
	assert RAM(12523) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(12523))))  severity failure;
	assert RAM(12524) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(12524))))  severity failure;
	assert RAM(12525) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(12525))))  severity failure;
	assert RAM(12526) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(12526))))  severity failure;
	assert RAM(12527) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(12527))))  severity failure;
	assert RAM(12528) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(12528))))  severity failure;
	assert RAM(12529) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(12529))))  severity failure;
	assert RAM(12530) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(12530))))  severity failure;
	assert RAM(12531) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(12531))))  severity failure;
	assert RAM(12532) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(12532))))  severity failure;
	assert RAM(12533) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(12533))))  severity failure;
	assert RAM(12534) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(12534))))  severity failure;
	assert RAM(12535) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(12535))))  severity failure;
	assert RAM(12536) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(12536))))  severity failure;
	assert RAM(12537) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(12537))))  severity failure;
	assert RAM(12538) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(12538))))  severity failure;
	assert RAM(12539) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(12539))))  severity failure;
	assert RAM(12540) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(12540))))  severity failure;
	assert RAM(12541) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(12541))))  severity failure;
	assert RAM(12542) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(12542))))  severity failure;
	assert RAM(12543) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(12543))))  severity failure;
	assert RAM(12544) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(12544))))  severity failure;
	assert RAM(12545) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(12545))))  severity failure;
	assert RAM(12546) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(12546))))  severity failure;
	assert RAM(12547) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(12547))))  severity failure;
	assert RAM(12548) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(12548))))  severity failure;
	assert RAM(12549) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(12549))))  severity failure;
	assert RAM(12550) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(12550))))  severity failure;
	assert RAM(12551) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(12551))))  severity failure;
	assert RAM(12552) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(12552))))  severity failure;
	assert RAM(12553) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(12553))))  severity failure;
	assert RAM(12554) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(12554))))  severity failure;
	assert RAM(12555) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(12555))))  severity failure;
	assert RAM(12556) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(12556))))  severity failure;
	assert RAM(12557) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(12557))))  severity failure;
	assert RAM(12558) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(12558))))  severity failure;
	assert RAM(12559) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(12559))))  severity failure;
	assert RAM(12560) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(12560))))  severity failure;
	assert RAM(12561) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(12561))))  severity failure;
	assert RAM(12562) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(12562))))  severity failure;
	assert RAM(12563) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(12563))))  severity failure;
	assert RAM(12564) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(12564))))  severity failure;
	assert RAM(12565) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(12565))))  severity failure;
	assert RAM(12566) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(12566))))  severity failure;
	assert RAM(12567) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(12567))))  severity failure;
	assert RAM(12568) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(12568))))  severity failure;
	assert RAM(12569) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(12569))))  severity failure;
	assert RAM(12570) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(12570))))  severity failure;
	assert RAM(12571) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(12571))))  severity failure;
	assert RAM(12572) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(12572))))  severity failure;
	assert RAM(12573) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(12573))))  severity failure;
	assert RAM(12574) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(12574))))  severity failure;
	assert RAM(12575) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(12575))))  severity failure;
	assert RAM(12576) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(12576))))  severity failure;
	assert RAM(12577) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(12577))))  severity failure;
	assert RAM(12578) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(12578))))  severity failure;
	assert RAM(12579) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(12579))))  severity failure;
	assert RAM(12580) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(12580))))  severity failure;
	assert RAM(12581) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(12581))))  severity failure;
	assert RAM(12582) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(12582))))  severity failure;
	assert RAM(12583) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(12583))))  severity failure;
	assert RAM(12584) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(12584))))  severity failure;
	assert RAM(12585) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(12585))))  severity failure;
	assert RAM(12586) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(12586))))  severity failure;
	assert RAM(12587) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(12587))))  severity failure;
	assert RAM(12588) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(12588))))  severity failure;
	assert RAM(12589) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(12589))))  severity failure;
	assert RAM(12590) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(12590))))  severity failure;
	assert RAM(12591) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(12591))))  severity failure;
	assert RAM(12592) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(12592))))  severity failure;
	assert RAM(12593) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(12593))))  severity failure;
	assert RAM(12594) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(12594))))  severity failure;
	assert RAM(12595) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(12595))))  severity failure;
	assert RAM(12596) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(12596))))  severity failure;
	assert RAM(12597) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(12597))))  severity failure;
	assert RAM(12598) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(12598))))  severity failure;
	assert RAM(12599) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(12599))))  severity failure;
	assert RAM(12600) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(12600))))  severity failure;
	assert RAM(12601) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(12601))))  severity failure;
	assert RAM(12602) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(12602))))  severity failure;
	assert RAM(12603) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(12603))))  severity failure;
	assert RAM(12604) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(12604))))  severity failure;
	assert RAM(12605) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(12605))))  severity failure;
	assert RAM(12606) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(12606))))  severity failure;
	assert RAM(12607) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(12607))))  severity failure;
	assert RAM(12608) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(12608))))  severity failure;
	assert RAM(12609) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(12609))))  severity failure;
	assert RAM(12610) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(12610))))  severity failure;
	assert RAM(12611) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(12611))))  severity failure;
	assert RAM(12612) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(12612))))  severity failure;
	assert RAM(12613) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(12613))))  severity failure;
	assert RAM(12614) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(12614))))  severity failure;
	assert RAM(12615) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(12615))))  severity failure;
	assert RAM(12616) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(12616))))  severity failure;
	assert RAM(12617) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(12617))))  severity failure;
	assert RAM(12618) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(12618))))  severity failure;
	assert RAM(12619) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(12619))))  severity failure;
	assert RAM(12620) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(12620))))  severity failure;
	assert RAM(12621) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(12621))))  severity failure;
	assert RAM(12622) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(12622))))  severity failure;
	assert RAM(12623) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(12623))))  severity failure;
	assert RAM(12624) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(12624))))  severity failure;
	assert RAM(12625) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(12625))))  severity failure;
	assert RAM(12626) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(12626))))  severity failure;
	assert RAM(12627) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(12627))))  severity failure;
	assert RAM(12628) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(12628))))  severity failure;
	assert RAM(12629) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(12629))))  severity failure;
	assert RAM(12630) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(12630))))  severity failure;
	assert RAM(12631) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(12631))))  severity failure;
	assert RAM(12632) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(12632))))  severity failure;
	assert RAM(12633) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(12633))))  severity failure;
	assert RAM(12634) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(12634))))  severity failure;
	assert RAM(12635) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(12635))))  severity failure;
	assert RAM(12636) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(12636))))  severity failure;
	assert RAM(12637) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(12637))))  severity failure;
	assert RAM(12638) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(12638))))  severity failure;
	assert RAM(12639) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(12639))))  severity failure;
	assert RAM(12640) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(12640))))  severity failure;
	assert RAM(12641) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(12641))))  severity failure;
	assert RAM(12642) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(12642))))  severity failure;
	assert RAM(12643) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(12643))))  severity failure;
	assert RAM(12644) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(12644))))  severity failure;
	assert RAM(12645) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(12645))))  severity failure;
	assert RAM(12646) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(12646))))  severity failure;
	assert RAM(12647) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(12647))))  severity failure;
	assert RAM(12648) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(12648))))  severity failure;
	assert RAM(12649) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(12649))))  severity failure;
	assert RAM(12650) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(12650))))  severity failure;
	assert RAM(12651) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(12651))))  severity failure;
	assert RAM(12652) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(12652))))  severity failure;
	assert RAM(12653) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(12653))))  severity failure;
	assert RAM(12654) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(12654))))  severity failure;
	assert RAM(12655) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(12655))))  severity failure;
	assert RAM(12656) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(12656))))  severity failure;
	assert RAM(12657) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(12657))))  severity failure;
	assert RAM(12658) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(12658))))  severity failure;
	assert RAM(12659) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(12659))))  severity failure;
	assert RAM(12660) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(12660))))  severity failure;
	assert RAM(12661) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(12661))))  severity failure;
	assert RAM(12662) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(12662))))  severity failure;
	assert RAM(12663) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(12663))))  severity failure;
	assert RAM(12664) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(12664))))  severity failure;
	assert RAM(12665) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(12665))))  severity failure;
	assert RAM(12666) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(12666))))  severity failure;
	assert RAM(12667) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(12667))))  severity failure;
	assert RAM(12668) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(12668))))  severity failure;
	assert RAM(12669) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(12669))))  severity failure;
	assert RAM(12670) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(12670))))  severity failure;
	assert RAM(12671) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(12671))))  severity failure;
	assert RAM(12672) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(12672))))  severity failure;
	assert RAM(12673) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(12673))))  severity failure;
	assert RAM(12674) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(12674))))  severity failure;
	assert RAM(12675) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(12675))))  severity failure;
	assert RAM(12676) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(12676))))  severity failure;
	assert RAM(12677) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(12677))))  severity failure;
	assert RAM(12678) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(12678))))  severity failure;
	assert RAM(12679) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(12679))))  severity failure;
	assert RAM(12680) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(12680))))  severity failure;
	assert RAM(12681) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(12681))))  severity failure;
	assert RAM(12682) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(12682))))  severity failure;
	assert RAM(12683) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(12683))))  severity failure;
	assert RAM(12684) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(12684))))  severity failure;
	assert RAM(12685) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(12685))))  severity failure;
	assert RAM(12686) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(12686))))  severity failure;
	assert RAM(12687) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(12687))))  severity failure;
	assert RAM(12688) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(12688))))  severity failure;
	assert RAM(12689) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(12689))))  severity failure;
	assert RAM(12690) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(12690))))  severity failure;
	assert RAM(12691) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(12691))))  severity failure;
	assert RAM(12692) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(12692))))  severity failure;
	assert RAM(12693) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(12693))))  severity failure;
	assert RAM(12694) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(12694))))  severity failure;
	assert RAM(12695) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(12695))))  severity failure;
	assert RAM(12696) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(12696))))  severity failure;
	assert RAM(12697) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(12697))))  severity failure;
	assert RAM(12698) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(12698))))  severity failure;
	assert RAM(12699) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(12699))))  severity failure;
	assert RAM(12700) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(12700))))  severity failure;
	assert RAM(12701) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(12701))))  severity failure;
	assert RAM(12702) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(12702))))  severity failure;
	assert RAM(12703) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(12703))))  severity failure;
	assert RAM(12704) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(12704))))  severity failure;
	assert RAM(12705) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(12705))))  severity failure;
	assert RAM(12706) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(12706))))  severity failure;
	assert RAM(12707) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(12707))))  severity failure;
	assert RAM(12708) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(12708))))  severity failure;
	assert RAM(12709) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(12709))))  severity failure;
	assert RAM(12710) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(12710))))  severity failure;
	assert RAM(12711) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(12711))))  severity failure;
	assert RAM(12712) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(12712))))  severity failure;
	assert RAM(12713) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(12713))))  severity failure;
	assert RAM(12714) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(12714))))  severity failure;
	assert RAM(12715) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(12715))))  severity failure;
	assert RAM(12716) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(12716))))  severity failure;
	assert RAM(12717) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(12717))))  severity failure;
	assert RAM(12718) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(12718))))  severity failure;
	assert RAM(12719) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(12719))))  severity failure;
	assert RAM(12720) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(12720))))  severity failure;
	assert RAM(12721) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(12721))))  severity failure;
	assert RAM(12722) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(12722))))  severity failure;
	assert RAM(12723) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(12723))))  severity failure;
	assert RAM(12724) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(12724))))  severity failure;
	assert RAM(12725) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(12725))))  severity failure;
	assert RAM(12726) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(12726))))  severity failure;
	assert RAM(12727) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(12727))))  severity failure;
	assert RAM(12728) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(12728))))  severity failure;
	assert RAM(12729) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(12729))))  severity failure;
	assert RAM(12730) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(12730))))  severity failure;
	assert RAM(12731) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(12731))))  severity failure;
	assert RAM(12732) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(12732))))  severity failure;
	assert RAM(12733) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(12733))))  severity failure;
	assert RAM(12734) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(12734))))  severity failure;
	assert RAM(12735) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(12735))))  severity failure;
	assert RAM(12736) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(12736))))  severity failure;
	assert RAM(12737) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(12737))))  severity failure;
	assert RAM(12738) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(12738))))  severity failure;
	assert RAM(12739) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(12739))))  severity failure;
	assert RAM(12740) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(12740))))  severity failure;
	assert RAM(12741) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(12741))))  severity failure;
	assert RAM(12742) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(12742))))  severity failure;
	assert RAM(12743) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(12743))))  severity failure;
	assert RAM(12744) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(12744))))  severity failure;
	assert RAM(12745) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(12745))))  severity failure;
	assert RAM(12746) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(12746))))  severity failure;
	assert RAM(12747) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(12747))))  severity failure;
	assert RAM(12748) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(12748))))  severity failure;
	assert RAM(12749) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(12749))))  severity failure;
	assert RAM(12750) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(12750))))  severity failure;
	assert RAM(12751) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(12751))))  severity failure;
	assert RAM(12752) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(12752))))  severity failure;
	assert RAM(12753) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(12753))))  severity failure;
	assert RAM(12754) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(12754))))  severity failure;
	assert RAM(12755) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(12755))))  severity failure;
	assert RAM(12756) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(12756))))  severity failure;
	assert RAM(12757) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(12757))))  severity failure;
	assert RAM(12758) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(12758))))  severity failure;
	assert RAM(12759) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(12759))))  severity failure;
	assert RAM(12760) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(12760))))  severity failure;
	assert RAM(12761) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(12761))))  severity failure;
	assert RAM(12762) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(12762))))  severity failure;
	assert RAM(12763) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(12763))))  severity failure;
	assert RAM(12764) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(12764))))  severity failure;
	assert RAM(12765) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(12765))))  severity failure;
	assert RAM(12766) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(12766))))  severity failure;
	assert RAM(12767) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(12767))))  severity failure;
	assert RAM(12768) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(12768))))  severity failure;
	assert RAM(12769) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(12769))))  severity failure;
	assert RAM(12770) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(12770))))  severity failure;
	assert RAM(12771) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(12771))))  severity failure;
	assert RAM(12772) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(12772))))  severity failure;
	assert RAM(12773) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(12773))))  severity failure;
	assert RAM(12774) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(12774))))  severity failure;
	assert RAM(12775) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(12775))))  severity failure;
	assert RAM(12776) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(12776))))  severity failure;
	assert RAM(12777) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(12777))))  severity failure;
	assert RAM(12778) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(12778))))  severity failure;
	assert RAM(12779) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(12779))))  severity failure;
	assert RAM(12780) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(12780))))  severity failure;
	assert RAM(12781) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(12781))))  severity failure;
	assert RAM(12782) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(12782))))  severity failure;
	assert RAM(12783) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(12783))))  severity failure;
	assert RAM(12784) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(12784))))  severity failure;
	assert RAM(12785) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(12785))))  severity failure;
	assert RAM(12786) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(12786))))  severity failure;
	assert RAM(12787) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(12787))))  severity failure;
	assert RAM(12788) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(12788))))  severity failure;
	assert RAM(12789) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(12789))))  severity failure;
	assert RAM(12790) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(12790))))  severity failure;
	assert RAM(12791) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(12791))))  severity failure;
	assert RAM(12792) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(12792))))  severity failure;
	assert RAM(12793) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(12793))))  severity failure;
	assert RAM(12794) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(12794))))  severity failure;
	assert RAM(12795) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(12795))))  severity failure;
	assert RAM(12796) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(12796))))  severity failure;
	assert RAM(12797) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(12797))))  severity failure;
	assert RAM(12798) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(12798))))  severity failure;
	assert RAM(12799) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(12799))))  severity failure;
	assert RAM(12800) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(12800))))  severity failure;
	assert RAM(12801) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(12801))))  severity failure;
	assert RAM(12802) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(12802))))  severity failure;
	assert RAM(12803) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(12803))))  severity failure;
	assert RAM(12804) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(12804))))  severity failure;
	assert RAM(12805) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(12805))))  severity failure;
	assert RAM(12806) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(12806))))  severity failure;
	assert RAM(12807) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(12807))))  severity failure;
	assert RAM(12808) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(12808))))  severity failure;
	assert RAM(12809) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(12809))))  severity failure;
	assert RAM(12810) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(12810))))  severity failure;
	assert RAM(12811) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(12811))))  severity failure;
	assert RAM(12812) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(12812))))  severity failure;
	assert RAM(12813) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(12813))))  severity failure;
	assert RAM(12814) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(12814))))  severity failure;
	assert RAM(12815) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(12815))))  severity failure;
	assert RAM(12816) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(12816))))  severity failure;
	assert RAM(12817) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(12817))))  severity failure;
	assert RAM(12818) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(12818))))  severity failure;
	assert RAM(12819) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(12819))))  severity failure;
	assert RAM(12820) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(12820))))  severity failure;
	assert RAM(12821) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(12821))))  severity failure;
	assert RAM(12822) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(12822))))  severity failure;
	assert RAM(12823) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(12823))))  severity failure;
	assert RAM(12824) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(12824))))  severity failure;
	assert RAM(12825) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(12825))))  severity failure;
	assert RAM(12826) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(12826))))  severity failure;
	assert RAM(12827) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(12827))))  severity failure;
	assert RAM(12828) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(12828))))  severity failure;
	assert RAM(12829) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(12829))))  severity failure;
	assert RAM(12830) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(12830))))  severity failure;
	assert RAM(12831) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(12831))))  severity failure;
	assert RAM(12832) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(12832))))  severity failure;
	assert RAM(12833) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(12833))))  severity failure;
	assert RAM(12834) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(12834))))  severity failure;
	assert RAM(12835) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(12835))))  severity failure;
	assert RAM(12836) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(12836))))  severity failure;
	assert RAM(12837) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(12837))))  severity failure;
	assert RAM(12838) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(12838))))  severity failure;
	assert RAM(12839) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(12839))))  severity failure;
	assert RAM(12840) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(12840))))  severity failure;
	assert RAM(12841) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(12841))))  severity failure;
	assert RAM(12842) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(12842))))  severity failure;
	assert RAM(12843) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(12843))))  severity failure;
	assert RAM(12844) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(12844))))  severity failure;
	assert RAM(12845) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(12845))))  severity failure;
	assert RAM(12846) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(12846))))  severity failure;
	assert RAM(12847) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(12847))))  severity failure;
	assert RAM(12848) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(12848))))  severity failure;
	assert RAM(12849) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(12849))))  severity failure;
	assert RAM(12850) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(12850))))  severity failure;
	assert RAM(12851) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(12851))))  severity failure;
	assert RAM(12852) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(12852))))  severity failure;
	assert RAM(12853) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(12853))))  severity failure;
	assert RAM(12854) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(12854))))  severity failure;
	assert RAM(12855) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(12855))))  severity failure;
	assert RAM(12856) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(12856))))  severity failure;
	assert RAM(12857) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(12857))))  severity failure;
	assert RAM(12858) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(12858))))  severity failure;
	assert RAM(12859) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(12859))))  severity failure;
	assert RAM(12860) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(12860))))  severity failure;
	assert RAM(12861) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(12861))))  severity failure;
	assert RAM(12862) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(12862))))  severity failure;
	assert RAM(12863) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(12863))))  severity failure;
	assert RAM(12864) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(12864))))  severity failure;
	assert RAM(12865) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(12865))))  severity failure;
	assert RAM(12866) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(12866))))  severity failure;
	assert RAM(12867) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(12867))))  severity failure;
	assert RAM(12868) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(12868))))  severity failure;
	assert RAM(12869) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(12869))))  severity failure;
	assert RAM(12870) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(12870))))  severity failure;
	assert RAM(12871) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(12871))))  severity failure;
	assert RAM(12872) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(12872))))  severity failure;
	assert RAM(12873) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(12873))))  severity failure;
	assert RAM(12874) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(12874))))  severity failure;
	assert RAM(12875) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(12875))))  severity failure;
	assert RAM(12876) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(12876))))  severity failure;
	assert RAM(12877) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(12877))))  severity failure;
	assert RAM(12878) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(12878))))  severity failure;
	assert RAM(12879) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(12879))))  severity failure;
	assert RAM(12880) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(12880))))  severity failure;
	assert RAM(12881) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(12881))))  severity failure;
	assert RAM(12882) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(12882))))  severity failure;
	assert RAM(12883) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(12883))))  severity failure;
	assert RAM(12884) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(12884))))  severity failure;
	assert RAM(12885) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(12885))))  severity failure;
	assert RAM(12886) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(12886))))  severity failure;
	assert RAM(12887) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(12887))))  severity failure;
	assert RAM(12888) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(12888))))  severity failure;
	assert RAM(12889) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(12889))))  severity failure;
	assert RAM(12890) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(12890))))  severity failure;
	assert RAM(12891) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(12891))))  severity failure;
	assert RAM(12892) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(12892))))  severity failure;
	assert RAM(12893) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(12893))))  severity failure;
	assert RAM(12894) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(12894))))  severity failure;
	assert RAM(12895) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(12895))))  severity failure;
	assert RAM(12896) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(12896))))  severity failure;
	assert RAM(12897) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(12897))))  severity failure;
	assert RAM(12898) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(12898))))  severity failure;
	assert RAM(12899) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(12899))))  severity failure;
	assert RAM(12900) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(12900))))  severity failure;
	assert RAM(12901) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(12901))))  severity failure;
	assert RAM(12902) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(12902))))  severity failure;
	assert RAM(12903) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(12903))))  severity failure;
	assert RAM(12904) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(12904))))  severity failure;
	assert RAM(12905) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(12905))))  severity failure;
	assert RAM(12906) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(12906))))  severity failure;
	assert RAM(12907) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(12907))))  severity failure;
	assert RAM(12908) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(12908))))  severity failure;
	assert RAM(12909) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(12909))))  severity failure;
	assert RAM(12910) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(12910))))  severity failure;
	assert RAM(12911) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(12911))))  severity failure;
	assert RAM(12912) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(12912))))  severity failure;
	assert RAM(12913) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(12913))))  severity failure;
	assert RAM(12914) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(12914))))  severity failure;
	assert RAM(12915) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(12915))))  severity failure;
	assert RAM(12916) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(12916))))  severity failure;
	assert RAM(12917) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(12917))))  severity failure;
	assert RAM(12918) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(12918))))  severity failure;
	assert RAM(12919) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(12919))))  severity failure;
	assert RAM(12920) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(12920))))  severity failure;
	assert RAM(12921) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(12921))))  severity failure;
	assert RAM(12922) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(12922))))  severity failure;
	assert RAM(12923) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(12923))))  severity failure;
	assert RAM(12924) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(12924))))  severity failure;
	assert RAM(12925) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(12925))))  severity failure;
	assert RAM(12926) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(12926))))  severity failure;
	assert RAM(12927) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(12927))))  severity failure;
	assert RAM(12928) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(12928))))  severity failure;
	assert RAM(12929) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(12929))))  severity failure;
	assert RAM(12930) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(12930))))  severity failure;
	assert RAM(12931) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(12931))))  severity failure;
	assert RAM(12932) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(12932))))  severity failure;
	assert RAM(12933) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(12933))))  severity failure;
	assert RAM(12934) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(12934))))  severity failure;
	assert RAM(12935) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(12935))))  severity failure;
	assert RAM(12936) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(12936))))  severity failure;
	assert RAM(12937) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(12937))))  severity failure;
	assert RAM(12938) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(12938))))  severity failure;
	assert RAM(12939) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(12939))))  severity failure;
	assert RAM(12940) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(12940))))  severity failure;
	assert RAM(12941) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(12941))))  severity failure;
	assert RAM(12942) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(12942))))  severity failure;
	assert RAM(12943) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(12943))))  severity failure;
	assert RAM(12944) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(12944))))  severity failure;
	assert RAM(12945) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(12945))))  severity failure;
	assert RAM(12946) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(12946))))  severity failure;
	assert RAM(12947) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(12947))))  severity failure;
	assert RAM(12948) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(12948))))  severity failure;
	assert RAM(12949) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(12949))))  severity failure;
	assert RAM(12950) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(12950))))  severity failure;
	assert RAM(12951) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(12951))))  severity failure;
	assert RAM(12952) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(12952))))  severity failure;
	assert RAM(12953) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(12953))))  severity failure;
	assert RAM(12954) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(12954))))  severity failure;
	assert RAM(12955) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(12955))))  severity failure;
	assert RAM(12956) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(12956))))  severity failure;
	assert RAM(12957) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(12957))))  severity failure;
	assert RAM(12958) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(12958))))  severity failure;
	assert RAM(12959) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(12959))))  severity failure;
	assert RAM(12960) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(12960))))  severity failure;
	assert RAM(12961) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(12961))))  severity failure;
	assert RAM(12962) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(12962))))  severity failure;
	assert RAM(12963) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(12963))))  severity failure;
	assert RAM(12964) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(12964))))  severity failure;
	assert RAM(12965) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(12965))))  severity failure;
	assert RAM(12966) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(12966))))  severity failure;
	assert RAM(12967) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(12967))))  severity failure;
	assert RAM(12968) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(12968))))  severity failure;
	assert RAM(12969) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(12969))))  severity failure;
	assert RAM(12970) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(12970))))  severity failure;
	assert RAM(12971) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(12971))))  severity failure;
	assert RAM(12972) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(12972))))  severity failure;
	assert RAM(12973) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(12973))))  severity failure;
	assert RAM(12974) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(12974))))  severity failure;
	assert RAM(12975) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(12975))))  severity failure;
	assert RAM(12976) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(12976))))  severity failure;
	assert RAM(12977) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(12977))))  severity failure;
	assert RAM(12978) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(12978))))  severity failure;
	assert RAM(12979) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(12979))))  severity failure;
	assert RAM(12980) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(12980))))  severity failure;
	assert RAM(12981) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(12981))))  severity failure;
	assert RAM(12982) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(12982))))  severity failure;
	assert RAM(12983) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(12983))))  severity failure;
	assert RAM(12984) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(12984))))  severity failure;
	assert RAM(12985) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(12985))))  severity failure;
	assert RAM(12986) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(12986))))  severity failure;
	assert RAM(12987) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(12987))))  severity failure;
	assert RAM(12988) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(12988))))  severity failure;
	assert RAM(12989) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(12989))))  severity failure;
	assert RAM(12990) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(12990))))  severity failure;
	assert RAM(12991) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(12991))))  severity failure;
	assert RAM(12992) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(12992))))  severity failure;
	assert RAM(12993) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(12993))))  severity failure;
	assert RAM(12994) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(12994))))  severity failure;
	assert RAM(12995) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(12995))))  severity failure;
	assert RAM(12996) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(12996))))  severity failure;
	assert RAM(12997) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(12997))))  severity failure;
	assert RAM(12998) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(12998))))  severity failure;
	assert RAM(12999) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(12999))))  severity failure;
	assert RAM(13000) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(13000))))  severity failure;
	assert RAM(13001) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(13001))))  severity failure;
	assert RAM(13002) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(13002))))  severity failure;
	assert RAM(13003) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(13003))))  severity failure;
	assert RAM(13004) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(13004))))  severity failure;
	assert RAM(13005) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(13005))))  severity failure;
	assert RAM(13006) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(13006))))  severity failure;
	assert RAM(13007) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(13007))))  severity failure;
	assert RAM(13008) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(13008))))  severity failure;
	assert RAM(13009) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(13009))))  severity failure;
	assert RAM(13010) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(13010))))  severity failure;
	assert RAM(13011) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(13011))))  severity failure;
	assert RAM(13012) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(13012))))  severity failure;
	assert RAM(13013) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(13013))))  severity failure;
	assert RAM(13014) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(13014))))  severity failure;
	assert RAM(13015) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(13015))))  severity failure;
	assert RAM(13016) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(13016))))  severity failure;
	assert RAM(13017) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(13017))))  severity failure;
	assert RAM(13018) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(13018))))  severity failure;
	assert RAM(13019) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(13019))))  severity failure;
	assert RAM(13020) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(13020))))  severity failure;
	assert RAM(13021) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(13021))))  severity failure;
	assert RAM(13022) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(13022))))  severity failure;
	assert RAM(13023) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(13023))))  severity failure;
	assert RAM(13024) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(13024))))  severity failure;
	assert RAM(13025) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(13025))))  severity failure;
	assert RAM(13026) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(13026))))  severity failure;
	assert RAM(13027) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(13027))))  severity failure;
	assert RAM(13028) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(13028))))  severity failure;
	assert RAM(13029) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(13029))))  severity failure;
	assert RAM(13030) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(13030))))  severity failure;
	assert RAM(13031) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(13031))))  severity failure;
	assert RAM(13032) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(13032))))  severity failure;
	assert RAM(13033) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(13033))))  severity failure;
	assert RAM(13034) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(13034))))  severity failure;
	assert RAM(13035) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(13035))))  severity failure;
	assert RAM(13036) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(13036))))  severity failure;
	assert RAM(13037) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(13037))))  severity failure;
	assert RAM(13038) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(13038))))  severity failure;
	assert RAM(13039) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(13039))))  severity failure;
	assert RAM(13040) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(13040))))  severity failure;
	assert RAM(13041) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(13041))))  severity failure;
	assert RAM(13042) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(13042))))  severity failure;
	assert RAM(13043) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(13043))))  severity failure;
	assert RAM(13044) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(13044))))  severity failure;
	assert RAM(13045) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(13045))))  severity failure;
	assert RAM(13046) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(13046))))  severity failure;
	assert RAM(13047) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(13047))))  severity failure;
	assert RAM(13048) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(13048))))  severity failure;
	assert RAM(13049) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(13049))))  severity failure;
	assert RAM(13050) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(13050))))  severity failure;
	assert RAM(13051) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(13051))))  severity failure;
	assert RAM(13052) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(13052))))  severity failure;
	assert RAM(13053) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(13053))))  severity failure;
	assert RAM(13054) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13054))))  severity failure;
	assert RAM(13055) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(13055))))  severity failure;
	assert RAM(13056) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(13056))))  severity failure;
	assert RAM(13057) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(13057))))  severity failure;
	assert RAM(13058) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(13058))))  severity failure;
	assert RAM(13059) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(13059))))  severity failure;
	assert RAM(13060) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(13060))))  severity failure;
	assert RAM(13061) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(13061))))  severity failure;
	assert RAM(13062) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(13062))))  severity failure;
	assert RAM(13063) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(13063))))  severity failure;
	assert RAM(13064) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(13064))))  severity failure;
	assert RAM(13065) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(13065))))  severity failure;
	assert RAM(13066) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(13066))))  severity failure;
	assert RAM(13067) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(13067))))  severity failure;
	assert RAM(13068) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(13068))))  severity failure;
	assert RAM(13069) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(13069))))  severity failure;
	assert RAM(13070) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(13070))))  severity failure;
	assert RAM(13071) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(13071))))  severity failure;
	assert RAM(13072) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(13072))))  severity failure;
	assert RAM(13073) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(13073))))  severity failure;
	assert RAM(13074) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(13074))))  severity failure;
	assert RAM(13075) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(13075))))  severity failure;
	assert RAM(13076) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(13076))))  severity failure;
	assert RAM(13077) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(13077))))  severity failure;
	assert RAM(13078) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(13078))))  severity failure;
	assert RAM(13079) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(13079))))  severity failure;
	assert RAM(13080) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(13080))))  severity failure;
	assert RAM(13081) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(13081))))  severity failure;
	assert RAM(13082) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(13082))))  severity failure;
	assert RAM(13083) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(13083))))  severity failure;
	assert RAM(13084) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(13084))))  severity failure;
	assert RAM(13085) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(13085))))  severity failure;
	assert RAM(13086) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(13086))))  severity failure;
	assert RAM(13087) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(13087))))  severity failure;
	assert RAM(13088) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(13088))))  severity failure;
	assert RAM(13089) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(13089))))  severity failure;
	assert RAM(13090) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(13090))))  severity failure;
	assert RAM(13091) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(13091))))  severity failure;
	assert RAM(13092) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(13092))))  severity failure;
	assert RAM(13093) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(13093))))  severity failure;
	assert RAM(13094) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(13094))))  severity failure;
	assert RAM(13095) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(13095))))  severity failure;
	assert RAM(13096) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(13096))))  severity failure;
	assert RAM(13097) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(13097))))  severity failure;
	assert RAM(13098) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(13098))))  severity failure;
	assert RAM(13099) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(13099))))  severity failure;
	assert RAM(13100) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(13100))))  severity failure;
	assert RAM(13101) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(13101))))  severity failure;
	assert RAM(13102) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(13102))))  severity failure;
	assert RAM(13103) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(13103))))  severity failure;
	assert RAM(13104) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(13104))))  severity failure;
	assert RAM(13105) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(13105))))  severity failure;
	assert RAM(13106) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(13106))))  severity failure;
	assert RAM(13107) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(13107))))  severity failure;
	assert RAM(13108) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(13108))))  severity failure;
	assert RAM(13109) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(13109))))  severity failure;
	assert RAM(13110) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(13110))))  severity failure;
	assert RAM(13111) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(13111))))  severity failure;
	assert RAM(13112) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(13112))))  severity failure;
	assert RAM(13113) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(13113))))  severity failure;
	assert RAM(13114) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(13114))))  severity failure;
	assert RAM(13115) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(13115))))  severity failure;
	assert RAM(13116) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(13116))))  severity failure;
	assert RAM(13117) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(13117))))  severity failure;
	assert RAM(13118) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(13118))))  severity failure;
	assert RAM(13119) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(13119))))  severity failure;
	assert RAM(13120) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(13120))))  severity failure;
	assert RAM(13121) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(13121))))  severity failure;
	assert RAM(13122) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(13122))))  severity failure;
	assert RAM(13123) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(13123))))  severity failure;
	assert RAM(13124) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(13124))))  severity failure;
	assert RAM(13125) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(13125))))  severity failure;
	assert RAM(13126) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(13126))))  severity failure;
	assert RAM(13127) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(13127))))  severity failure;
	assert RAM(13128) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(13128))))  severity failure;
	assert RAM(13129) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(13129))))  severity failure;
	assert RAM(13130) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(13130))))  severity failure;
	assert RAM(13131) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(13131))))  severity failure;
	assert RAM(13132) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(13132))))  severity failure;
	assert RAM(13133) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(13133))))  severity failure;
	assert RAM(13134) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(13134))))  severity failure;
	assert RAM(13135) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(13135))))  severity failure;
	assert RAM(13136) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(13136))))  severity failure;
	assert RAM(13137) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(13137))))  severity failure;
	assert RAM(13138) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(13138))))  severity failure;
	assert RAM(13139) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(13139))))  severity failure;
	assert RAM(13140) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(13140))))  severity failure;
	assert RAM(13141) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(13141))))  severity failure;
	assert RAM(13142) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(13142))))  severity failure;
	assert RAM(13143) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(13143))))  severity failure;
	assert RAM(13144) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(13144))))  severity failure;
	assert RAM(13145) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(13145))))  severity failure;
	assert RAM(13146) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13146))))  severity failure;
	assert RAM(13147) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(13147))))  severity failure;
	assert RAM(13148) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(13148))))  severity failure;
	assert RAM(13149) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(13149))))  severity failure;
	assert RAM(13150) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(13150))))  severity failure;
	assert RAM(13151) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(13151))))  severity failure;
	assert RAM(13152) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(13152))))  severity failure;
	assert RAM(13153) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(13153))))  severity failure;
	assert RAM(13154) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(13154))))  severity failure;
	assert RAM(13155) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(13155))))  severity failure;
	assert RAM(13156) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(13156))))  severity failure;
	assert RAM(13157) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(13157))))  severity failure;
	assert RAM(13158) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(13158))))  severity failure;
	assert RAM(13159) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(13159))))  severity failure;
	assert RAM(13160) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(13160))))  severity failure;
	assert RAM(13161) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(13161))))  severity failure;
	assert RAM(13162) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(13162))))  severity failure;
	assert RAM(13163) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(13163))))  severity failure;
	assert RAM(13164) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(13164))))  severity failure;
	assert RAM(13165) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(13165))))  severity failure;
	assert RAM(13166) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(13166))))  severity failure;
	assert RAM(13167) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(13167))))  severity failure;
	assert RAM(13168) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(13168))))  severity failure;
	assert RAM(13169) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(13169))))  severity failure;
	assert RAM(13170) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(13170))))  severity failure;
	assert RAM(13171) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(13171))))  severity failure;
	assert RAM(13172) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(13172))))  severity failure;
	assert RAM(13173) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(13173))))  severity failure;
	assert RAM(13174) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(13174))))  severity failure;
	assert RAM(13175) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(13175))))  severity failure;
	assert RAM(13176) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(13176))))  severity failure;
	assert RAM(13177) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(13177))))  severity failure;
	assert RAM(13178) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(13178))))  severity failure;
	assert RAM(13179) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(13179))))  severity failure;
	assert RAM(13180) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(13180))))  severity failure;
	assert RAM(13181) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(13181))))  severity failure;
	assert RAM(13182) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(13182))))  severity failure;
	assert RAM(13183) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(13183))))  severity failure;
	assert RAM(13184) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(13184))))  severity failure;
	assert RAM(13185) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(13185))))  severity failure;
	assert RAM(13186) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(13186))))  severity failure;
	assert RAM(13187) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(13187))))  severity failure;
	assert RAM(13188) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(13188))))  severity failure;
	assert RAM(13189) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(13189))))  severity failure;
	assert RAM(13190) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(13190))))  severity failure;
	assert RAM(13191) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(13191))))  severity failure;
	assert RAM(13192) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(13192))))  severity failure;
	assert RAM(13193) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(13193))))  severity failure;
	assert RAM(13194) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(13194))))  severity failure;
	assert RAM(13195) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(13195))))  severity failure;
	assert RAM(13196) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(13196))))  severity failure;
	assert RAM(13197) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(13197))))  severity failure;
	assert RAM(13198) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(13198))))  severity failure;
	assert RAM(13199) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(13199))))  severity failure;
	assert RAM(13200) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(13200))))  severity failure;
	assert RAM(13201) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(13201))))  severity failure;
	assert RAM(13202) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(13202))))  severity failure;
	assert RAM(13203) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(13203))))  severity failure;
	assert RAM(13204) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(13204))))  severity failure;
	assert RAM(13205) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(13205))))  severity failure;
	assert RAM(13206) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(13206))))  severity failure;
	assert RAM(13207) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(13207))))  severity failure;
	assert RAM(13208) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(13208))))  severity failure;
	assert RAM(13209) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(13209))))  severity failure;
	assert RAM(13210) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(13210))))  severity failure;
	assert RAM(13211) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(13211))))  severity failure;
	assert RAM(13212) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(13212))))  severity failure;
	assert RAM(13213) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(13213))))  severity failure;
	assert RAM(13214) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(13214))))  severity failure;
	assert RAM(13215) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(13215))))  severity failure;
	assert RAM(13216) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(13216))))  severity failure;
	assert RAM(13217) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(13217))))  severity failure;
	assert RAM(13218) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(13218))))  severity failure;
	assert RAM(13219) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(13219))))  severity failure;
	assert RAM(13220) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(13220))))  severity failure;
	assert RAM(13221) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(13221))))  severity failure;
	assert RAM(13222) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(13222))))  severity failure;
	assert RAM(13223) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(13223))))  severity failure;
	assert RAM(13224) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(13224))))  severity failure;
	assert RAM(13225) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(13225))))  severity failure;
	assert RAM(13226) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(13226))))  severity failure;
	assert RAM(13227) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(13227))))  severity failure;
	assert RAM(13228) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(13228))))  severity failure;
	assert RAM(13229) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13229))))  severity failure;
	assert RAM(13230) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(13230))))  severity failure;
	assert RAM(13231) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(13231))))  severity failure;
	assert RAM(13232) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(13232))))  severity failure;
	assert RAM(13233) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(13233))))  severity failure;
	assert RAM(13234) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(13234))))  severity failure;
	assert RAM(13235) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(13235))))  severity failure;
	assert RAM(13236) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(13236))))  severity failure;
	assert RAM(13237) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(13237))))  severity failure;
	assert RAM(13238) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(13238))))  severity failure;
	assert RAM(13239) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(13239))))  severity failure;
	assert RAM(13240) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(13240))))  severity failure;
	assert RAM(13241) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(13241))))  severity failure;
	assert RAM(13242) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(13242))))  severity failure;
	assert RAM(13243) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(13243))))  severity failure;
	assert RAM(13244) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(13244))))  severity failure;
	assert RAM(13245) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(13245))))  severity failure;
	assert RAM(13246) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(13246))))  severity failure;
	assert RAM(13247) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(13247))))  severity failure;
	assert RAM(13248) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(13248))))  severity failure;
	assert RAM(13249) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(13249))))  severity failure;
	assert RAM(13250) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(13250))))  severity failure;
	assert RAM(13251) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(13251))))  severity failure;
	assert RAM(13252) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(13252))))  severity failure;
	assert RAM(13253) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(13253))))  severity failure;
	assert RAM(13254) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(13254))))  severity failure;
	assert RAM(13255) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(13255))))  severity failure;
	assert RAM(13256) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(13256))))  severity failure;
	assert RAM(13257) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(13257))))  severity failure;
	assert RAM(13258) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(13258))))  severity failure;
	assert RAM(13259) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(13259))))  severity failure;
	assert RAM(13260) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(13260))))  severity failure;
	assert RAM(13261) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(13261))))  severity failure;
	assert RAM(13262) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(13262))))  severity failure;
	assert RAM(13263) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(13263))))  severity failure;
	assert RAM(13264) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(13264))))  severity failure;
	assert RAM(13265) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(13265))))  severity failure;
	assert RAM(13266) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(13266))))  severity failure;
	assert RAM(13267) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(13267))))  severity failure;
	assert RAM(13268) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(13268))))  severity failure;
	assert RAM(13269) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(13269))))  severity failure;
	assert RAM(13270) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(13270))))  severity failure;
	assert RAM(13271) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(13271))))  severity failure;
	assert RAM(13272) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(13272))))  severity failure;
	assert RAM(13273) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(13273))))  severity failure;
	assert RAM(13274) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(13274))))  severity failure;
	assert RAM(13275) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(13275))))  severity failure;
	assert RAM(13276) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(13276))))  severity failure;
	assert RAM(13277) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(13277))))  severity failure;
	assert RAM(13278) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(13278))))  severity failure;
	assert RAM(13279) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(13279))))  severity failure;
	assert RAM(13280) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(13280))))  severity failure;
	assert RAM(13281) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(13281))))  severity failure;
	assert RAM(13282) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(13282))))  severity failure;
	assert RAM(13283) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(13283))))  severity failure;
	assert RAM(13284) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(13284))))  severity failure;
	assert RAM(13285) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(13285))))  severity failure;
	assert RAM(13286) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(13286))))  severity failure;
	assert RAM(13287) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(13287))))  severity failure;
	assert RAM(13288) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(13288))))  severity failure;
	assert RAM(13289) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(13289))))  severity failure;
	assert RAM(13290) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(13290))))  severity failure;
	assert RAM(13291) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(13291))))  severity failure;
	assert RAM(13292) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(13292))))  severity failure;
	assert RAM(13293) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(13293))))  severity failure;
	assert RAM(13294) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(13294))))  severity failure;
	assert RAM(13295) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(13295))))  severity failure;
	assert RAM(13296) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(13296))))  severity failure;
	assert RAM(13297) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(13297))))  severity failure;
	assert RAM(13298) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(13298))))  severity failure;
	assert RAM(13299) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(13299))))  severity failure;
	assert RAM(13300) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(13300))))  severity failure;
	assert RAM(13301) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(13301))))  severity failure;
	assert RAM(13302) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(13302))))  severity failure;
	assert RAM(13303) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(13303))))  severity failure;
	assert RAM(13304) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(13304))))  severity failure;
	assert RAM(13305) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(13305))))  severity failure;
	assert RAM(13306) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(13306))))  severity failure;
	assert RAM(13307) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(13307))))  severity failure;
	assert RAM(13308) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(13308))))  severity failure;
	assert RAM(13309) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(13309))))  severity failure;
	assert RAM(13310) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(13310))))  severity failure;
	assert RAM(13311) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(13311))))  severity failure;
	assert RAM(13312) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(13312))))  severity failure;
	assert RAM(13313) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(13313))))  severity failure;
	assert RAM(13314) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(13314))))  severity failure;
	assert RAM(13315) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(13315))))  severity failure;
	assert RAM(13316) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(13316))))  severity failure;
	assert RAM(13317) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(13317))))  severity failure;
	assert RAM(13318) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(13318))))  severity failure;
	assert RAM(13319) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(13319))))  severity failure;
	assert RAM(13320) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(13320))))  severity failure;
	assert RAM(13321) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(13321))))  severity failure;
	assert RAM(13322) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(13322))))  severity failure;
	assert RAM(13323) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(13323))))  severity failure;
	assert RAM(13324) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(13324))))  severity failure;
	assert RAM(13325) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(13325))))  severity failure;
	assert RAM(13326) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(13326))))  severity failure;
	assert RAM(13327) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(13327))))  severity failure;
	assert RAM(13328) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(13328))))  severity failure;
	assert RAM(13329) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(13329))))  severity failure;
	assert RAM(13330) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(13330))))  severity failure;
	assert RAM(13331) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(13331))))  severity failure;
	assert RAM(13332) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(13332))))  severity failure;
	assert RAM(13333) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(13333))))  severity failure;
	assert RAM(13334) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(13334))))  severity failure;
	assert RAM(13335) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(13335))))  severity failure;
	assert RAM(13336) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(13336))))  severity failure;
	assert RAM(13337) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(13337))))  severity failure;
	assert RAM(13338) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(13338))))  severity failure;
	assert RAM(13339) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(13339))))  severity failure;
	assert RAM(13340) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(13340))))  severity failure;
	assert RAM(13341) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(13341))))  severity failure;
	assert RAM(13342) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(13342))))  severity failure;
	assert RAM(13343) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(13343))))  severity failure;
	assert RAM(13344) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(13344))))  severity failure;
	assert RAM(13345) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(13345))))  severity failure;
	assert RAM(13346) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(13346))))  severity failure;
	assert RAM(13347) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(13347))))  severity failure;
	assert RAM(13348) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(13348))))  severity failure;
	assert RAM(13349) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(13349))))  severity failure;
	assert RAM(13350) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(13350))))  severity failure;
	assert RAM(13351) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(13351))))  severity failure;
	assert RAM(13352) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(13352))))  severity failure;
	assert RAM(13353) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(13353))))  severity failure;
	assert RAM(13354) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(13354))))  severity failure;
	assert RAM(13355) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(13355))))  severity failure;
	assert RAM(13356) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(13356))))  severity failure;
	assert RAM(13357) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(13357))))  severity failure;
	assert RAM(13358) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(13358))))  severity failure;
	assert RAM(13359) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(13359))))  severity failure;
	assert RAM(13360) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(13360))))  severity failure;
	assert RAM(13361) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(13361))))  severity failure;
	assert RAM(13362) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(13362))))  severity failure;
	assert RAM(13363) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(13363))))  severity failure;
	assert RAM(13364) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(13364))))  severity failure;
	assert RAM(13365) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(13365))))  severity failure;
	assert RAM(13366) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(13366))))  severity failure;
	assert RAM(13367) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(13367))))  severity failure;
	assert RAM(13368) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(13368))))  severity failure;
	assert RAM(13369) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(13369))))  severity failure;
	assert RAM(13370) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(13370))))  severity failure;
	assert RAM(13371) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(13371))))  severity failure;
	assert RAM(13372) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(13372))))  severity failure;
	assert RAM(13373) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(13373))))  severity failure;
	assert RAM(13374) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(13374))))  severity failure;
	assert RAM(13375) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(13375))))  severity failure;
	assert RAM(13376) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(13376))))  severity failure;
	assert RAM(13377) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(13377))))  severity failure;
	assert RAM(13378) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(13378))))  severity failure;
	assert RAM(13379) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(13379))))  severity failure;
	assert RAM(13380) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(13380))))  severity failure;
	assert RAM(13381) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(13381))))  severity failure;
	assert RAM(13382) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(13382))))  severity failure;
	assert RAM(13383) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(13383))))  severity failure;
	assert RAM(13384) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(13384))))  severity failure;
	assert RAM(13385) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(13385))))  severity failure;
	assert RAM(13386) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(13386))))  severity failure;
	assert RAM(13387) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(13387))))  severity failure;
	assert RAM(13388) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(13388))))  severity failure;
	assert RAM(13389) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(13389))))  severity failure;
	assert RAM(13390) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(13390))))  severity failure;
	assert RAM(13391) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(13391))))  severity failure;
	assert RAM(13392) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(13392))))  severity failure;
	assert RAM(13393) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(13393))))  severity failure;
	assert RAM(13394) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(13394))))  severity failure;
	assert RAM(13395) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(13395))))  severity failure;
	assert RAM(13396) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(13396))))  severity failure;
	assert RAM(13397) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(13397))))  severity failure;
	assert RAM(13398) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(13398))))  severity failure;
	assert RAM(13399) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(13399))))  severity failure;
	assert RAM(13400) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(13400))))  severity failure;
	assert RAM(13401) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(13401))))  severity failure;
	assert RAM(13402) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(13402))))  severity failure;
	assert RAM(13403) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(13403))))  severity failure;
	assert RAM(13404) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(13404))))  severity failure;
	assert RAM(13405) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(13405))))  severity failure;
	assert RAM(13406) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(13406))))  severity failure;
	assert RAM(13407) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(13407))))  severity failure;
	assert RAM(13408) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(13408))))  severity failure;
	assert RAM(13409) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(13409))))  severity failure;
	assert RAM(13410) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(13410))))  severity failure;
	assert RAM(13411) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(13411))))  severity failure;
	assert RAM(13412) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(13412))))  severity failure;
	assert RAM(13413) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(13413))))  severity failure;
	assert RAM(13414) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(13414))))  severity failure;
	assert RAM(13415) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(13415))))  severity failure;
	assert RAM(13416) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(13416))))  severity failure;
	assert RAM(13417) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(13417))))  severity failure;
	assert RAM(13418) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(13418))))  severity failure;
	assert RAM(13419) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(13419))))  severity failure;
	assert RAM(13420) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(13420))))  severity failure;
	assert RAM(13421) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(13421))))  severity failure;
	assert RAM(13422) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(13422))))  severity failure;
	assert RAM(13423) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(13423))))  severity failure;
	assert RAM(13424) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(13424))))  severity failure;
	assert RAM(13425) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13425))))  severity failure;
	assert RAM(13426) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(13426))))  severity failure;
	assert RAM(13427) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(13427))))  severity failure;
	assert RAM(13428) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(13428))))  severity failure;
	assert RAM(13429) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(13429))))  severity failure;
	assert RAM(13430) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(13430))))  severity failure;
	assert RAM(13431) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(13431))))  severity failure;
	assert RAM(13432) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(13432))))  severity failure;
	assert RAM(13433) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(13433))))  severity failure;
	assert RAM(13434) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(13434))))  severity failure;
	assert RAM(13435) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(13435))))  severity failure;
	assert RAM(13436) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(13436))))  severity failure;
	assert RAM(13437) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(13437))))  severity failure;
	assert RAM(13438) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(13438))))  severity failure;
	assert RAM(13439) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(13439))))  severity failure;
	assert RAM(13440) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(13440))))  severity failure;
	assert RAM(13441) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(13441))))  severity failure;
	assert RAM(13442) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(13442))))  severity failure;
	assert RAM(13443) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(13443))))  severity failure;
	assert RAM(13444) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(13444))))  severity failure;
	assert RAM(13445) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(13445))))  severity failure;
	assert RAM(13446) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(13446))))  severity failure;
	assert RAM(13447) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13447))))  severity failure;
	assert RAM(13448) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(13448))))  severity failure;
	assert RAM(13449) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(13449))))  severity failure;
	assert RAM(13450) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(13450))))  severity failure;
	assert RAM(13451) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(13451))))  severity failure;
	assert RAM(13452) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(13452))))  severity failure;
	assert RAM(13453) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(13453))))  severity failure;
	assert RAM(13454) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(13454))))  severity failure;
	assert RAM(13455) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(13455))))  severity failure;
	assert RAM(13456) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(13456))))  severity failure;
	assert RAM(13457) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(13457))))  severity failure;
	assert RAM(13458) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(13458))))  severity failure;
	assert RAM(13459) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(13459))))  severity failure;
	assert RAM(13460) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(13460))))  severity failure;
	assert RAM(13461) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(13461))))  severity failure;
	assert RAM(13462) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(13462))))  severity failure;
	assert RAM(13463) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(13463))))  severity failure;
	assert RAM(13464) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(13464))))  severity failure;
	assert RAM(13465) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(13465))))  severity failure;
	assert RAM(13466) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(13466))))  severity failure;
	assert RAM(13467) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(13467))))  severity failure;
	assert RAM(13468) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(13468))))  severity failure;
	assert RAM(13469) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(13469))))  severity failure;
	assert RAM(13470) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(13470))))  severity failure;
	assert RAM(13471) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(13471))))  severity failure;
	assert RAM(13472) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(13472))))  severity failure;
	assert RAM(13473) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(13473))))  severity failure;
	assert RAM(13474) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(13474))))  severity failure;
	assert RAM(13475) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(13475))))  severity failure;
	assert RAM(13476) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(13476))))  severity failure;
	assert RAM(13477) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(13477))))  severity failure;
	assert RAM(13478) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(13478))))  severity failure;
	assert RAM(13479) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(13479))))  severity failure;
	assert RAM(13480) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(13480))))  severity failure;
	assert RAM(13481) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(13481))))  severity failure;
	assert RAM(13482) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(13482))))  severity failure;
	assert RAM(13483) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(13483))))  severity failure;
	assert RAM(13484) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(13484))))  severity failure;
	assert RAM(13485) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(13485))))  severity failure;
	assert RAM(13486) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(13486))))  severity failure;
	assert RAM(13487) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(13487))))  severity failure;
	assert RAM(13488) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(13488))))  severity failure;
	assert RAM(13489) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(13489))))  severity failure;
	assert RAM(13490) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(13490))))  severity failure;
	assert RAM(13491) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(13491))))  severity failure;
	assert RAM(13492) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(13492))))  severity failure;
	assert RAM(13493) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(13493))))  severity failure;
	assert RAM(13494) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(13494))))  severity failure;
	assert RAM(13495) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(13495))))  severity failure;
	assert RAM(13496) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(13496))))  severity failure;
	assert RAM(13497) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(13497))))  severity failure;
	assert RAM(13498) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(13498))))  severity failure;
	assert RAM(13499) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(13499))))  severity failure;
	assert RAM(13500) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(13500))))  severity failure;
	assert RAM(13501) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(13501))))  severity failure;
	assert RAM(13502) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(13502))))  severity failure;
	assert RAM(13503) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(13503))))  severity failure;
	assert RAM(13504) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(13504))))  severity failure;
	assert RAM(13505) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(13505))))  severity failure;
	assert RAM(13506) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(13506))))  severity failure;
	assert RAM(13507) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(13507))))  severity failure;
	assert RAM(13508) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(13508))))  severity failure;
	assert RAM(13509) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(13509))))  severity failure;
	assert RAM(13510) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(13510))))  severity failure;
	assert RAM(13511) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(13511))))  severity failure;
	assert RAM(13512) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(13512))))  severity failure;
	assert RAM(13513) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(13513))))  severity failure;
	assert RAM(13514) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(13514))))  severity failure;
	assert RAM(13515) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(13515))))  severity failure;
	assert RAM(13516) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(13516))))  severity failure;
	assert RAM(13517) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(13517))))  severity failure;
	assert RAM(13518) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(13518))))  severity failure;
	assert RAM(13519) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(13519))))  severity failure;
	assert RAM(13520) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(13520))))  severity failure;
	assert RAM(13521) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(13521))))  severity failure;
	assert RAM(13522) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(13522))))  severity failure;
	assert RAM(13523) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(13523))))  severity failure;
	assert RAM(13524) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(13524))))  severity failure;
	assert RAM(13525) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(13525))))  severity failure;
	assert RAM(13526) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(13526))))  severity failure;
	assert RAM(13527) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(13527))))  severity failure;
	assert RAM(13528) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(13528))))  severity failure;
	assert RAM(13529) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(13529))))  severity failure;
	assert RAM(13530) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(13530))))  severity failure;
	assert RAM(13531) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(13531))))  severity failure;
	assert RAM(13532) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(13532))))  severity failure;
	assert RAM(13533) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(13533))))  severity failure;
	assert RAM(13534) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(13534))))  severity failure;
	assert RAM(13535) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(13535))))  severity failure;
	assert RAM(13536) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(13536))))  severity failure;
	assert RAM(13537) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(13537))))  severity failure;
	assert RAM(13538) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(13538))))  severity failure;
	assert RAM(13539) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(13539))))  severity failure;
	assert RAM(13540) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(13540))))  severity failure;
	assert RAM(13541) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(13541))))  severity failure;
	assert RAM(13542) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(13542))))  severity failure;
	assert RAM(13543) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(13543))))  severity failure;
	assert RAM(13544) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(13544))))  severity failure;
	assert RAM(13545) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(13545))))  severity failure;
	assert RAM(13546) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(13546))))  severity failure;
	assert RAM(13547) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(13547))))  severity failure;
	assert RAM(13548) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(13548))))  severity failure;
	assert RAM(13549) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(13549))))  severity failure;
	assert RAM(13550) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(13550))))  severity failure;
	assert RAM(13551) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(13551))))  severity failure;
	assert RAM(13552) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(13552))))  severity failure;
	assert RAM(13553) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(13553))))  severity failure;
	assert RAM(13554) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(13554))))  severity failure;
	assert RAM(13555) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(13555))))  severity failure;
	assert RAM(13556) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(13556))))  severity failure;
	assert RAM(13557) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(13557))))  severity failure;
	assert RAM(13558) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(13558))))  severity failure;
	assert RAM(13559) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(13559))))  severity failure;
	assert RAM(13560) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(13560))))  severity failure;
	assert RAM(13561) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(13561))))  severity failure;
	assert RAM(13562) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(13562))))  severity failure;
	assert RAM(13563) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(13563))))  severity failure;
	assert RAM(13564) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(13564))))  severity failure;
	assert RAM(13565) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(13565))))  severity failure;
	assert RAM(13566) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(13566))))  severity failure;
	assert RAM(13567) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(13567))))  severity failure;
	assert RAM(13568) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(13568))))  severity failure;
	assert RAM(13569) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(13569))))  severity failure;
	assert RAM(13570) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(13570))))  severity failure;
	assert RAM(13571) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(13571))))  severity failure;
	assert RAM(13572) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(13572))))  severity failure;
	assert RAM(13573) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(13573))))  severity failure;
	assert RAM(13574) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(13574))))  severity failure;
	assert RAM(13575) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(13575))))  severity failure;
	assert RAM(13576) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(13576))))  severity failure;
	assert RAM(13577) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(13577))))  severity failure;
	assert RAM(13578) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(13578))))  severity failure;
	assert RAM(13579) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(13579))))  severity failure;
	assert RAM(13580) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(13580))))  severity failure;
	assert RAM(13581) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(13581))))  severity failure;
	assert RAM(13582) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(13582))))  severity failure;
	assert RAM(13583) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(13583))))  severity failure;
	assert RAM(13584) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(13584))))  severity failure;
	assert RAM(13585) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(13585))))  severity failure;
	assert RAM(13586) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(13586))))  severity failure;
	assert RAM(13587) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(13587))))  severity failure;
	assert RAM(13588) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(13588))))  severity failure;
	assert RAM(13589) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(13589))))  severity failure;
	assert RAM(13590) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(13590))))  severity failure;
	assert RAM(13591) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(13591))))  severity failure;
	assert RAM(13592) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(13592))))  severity failure;
	assert RAM(13593) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(13593))))  severity failure;
	assert RAM(13594) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(13594))))  severity failure;
	assert RAM(13595) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(13595))))  severity failure;
	assert RAM(13596) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(13596))))  severity failure;
	assert RAM(13597) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(13597))))  severity failure;
	assert RAM(13598) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(13598))))  severity failure;
	assert RAM(13599) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(13599))))  severity failure;
	assert RAM(13600) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(13600))))  severity failure;
	assert RAM(13601) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(13601))))  severity failure;
	assert RAM(13602) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(13602))))  severity failure;
	assert RAM(13603) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(13603))))  severity failure;
	assert RAM(13604) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(13604))))  severity failure;
	assert RAM(13605) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(13605))))  severity failure;
	assert RAM(13606) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(13606))))  severity failure;
	assert RAM(13607) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(13607))))  severity failure;
	assert RAM(13608) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(13608))))  severity failure;
	assert RAM(13609) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(13609))))  severity failure;
	assert RAM(13610) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(13610))))  severity failure;
	assert RAM(13611) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(13611))))  severity failure;
	assert RAM(13612) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(13612))))  severity failure;
	assert RAM(13613) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(13613))))  severity failure;
	assert RAM(13614) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(13614))))  severity failure;
	assert RAM(13615) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(13615))))  severity failure;
	assert RAM(13616) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(13616))))  severity failure;
	assert RAM(13617) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(13617))))  severity failure;
	assert RAM(13618) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(13618))))  severity failure;
	assert RAM(13619) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(13619))))  severity failure;
	assert RAM(13620) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(13620))))  severity failure;
	assert RAM(13621) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(13621))))  severity failure;
	assert RAM(13622) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(13622))))  severity failure;
	assert RAM(13623) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(13623))))  severity failure;
	assert RAM(13624) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(13624))))  severity failure;
	assert RAM(13625) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(13625))))  severity failure;
	assert RAM(13626) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(13626))))  severity failure;
	assert RAM(13627) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(13627))))  severity failure;
	assert RAM(13628) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(13628))))  severity failure;
	assert RAM(13629) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(13629))))  severity failure;
	assert RAM(13630) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(13630))))  severity failure;
	assert RAM(13631) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(13631))))  severity failure;
	assert RAM(13632) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(13632))))  severity failure;
	assert RAM(13633) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(13633))))  severity failure;
	assert RAM(13634) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(13634))))  severity failure;
	assert RAM(13635) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(13635))))  severity failure;
	assert RAM(13636) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(13636))))  severity failure;
	assert RAM(13637) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(13637))))  severity failure;
	assert RAM(13638) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(13638))))  severity failure;
	assert RAM(13639) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(13639))))  severity failure;
	assert RAM(13640) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(13640))))  severity failure;
	assert RAM(13641) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(13641))))  severity failure;
	assert RAM(13642) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(13642))))  severity failure;
	assert RAM(13643) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(13643))))  severity failure;
	assert RAM(13644) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(13644))))  severity failure;
	assert RAM(13645) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(13645))))  severity failure;
	assert RAM(13646) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(13646))))  severity failure;
	assert RAM(13647) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(13647))))  severity failure;
	assert RAM(13648) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(13648))))  severity failure;
	assert RAM(13649) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(13649))))  severity failure;
	assert RAM(13650) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(13650))))  severity failure;
	assert RAM(13651) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(13651))))  severity failure;
	assert RAM(13652) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(13652))))  severity failure;
	assert RAM(13653) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(13653))))  severity failure;
	assert RAM(13654) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(13654))))  severity failure;
	assert RAM(13655) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(13655))))  severity failure;
	assert RAM(13656) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(13656))))  severity failure;
	assert RAM(13657) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(13657))))  severity failure;
	assert RAM(13658) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(13658))))  severity failure;
	assert RAM(13659) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(13659))))  severity failure;
	assert RAM(13660) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(13660))))  severity failure;
	assert RAM(13661) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(13661))))  severity failure;
	assert RAM(13662) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(13662))))  severity failure;
	assert RAM(13663) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(13663))))  severity failure;
	assert RAM(13664) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(13664))))  severity failure;
	assert RAM(13665) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(13665))))  severity failure;
	assert RAM(13666) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(13666))))  severity failure;
	assert RAM(13667) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(13667))))  severity failure;
	assert RAM(13668) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(13668))))  severity failure;
	assert RAM(13669) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(13669))))  severity failure;
	assert RAM(13670) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(13670))))  severity failure;
	assert RAM(13671) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(13671))))  severity failure;
	assert RAM(13672) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(13672))))  severity failure;
	assert RAM(13673) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(13673))))  severity failure;
	assert RAM(13674) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(13674))))  severity failure;
	assert RAM(13675) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(13675))))  severity failure;
	assert RAM(13676) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(13676))))  severity failure;
	assert RAM(13677) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(13677))))  severity failure;
	assert RAM(13678) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(13678))))  severity failure;
	assert RAM(13679) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(13679))))  severity failure;
	assert RAM(13680) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(13680))))  severity failure;
	assert RAM(13681) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(13681))))  severity failure;
	assert RAM(13682) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(13682))))  severity failure;
	assert RAM(13683) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(13683))))  severity failure;
	assert RAM(13684) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(13684))))  severity failure;
	assert RAM(13685) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(13685))))  severity failure;
	assert RAM(13686) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(13686))))  severity failure;
	assert RAM(13687) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(13687))))  severity failure;
	assert RAM(13688) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(13688))))  severity failure;
	assert RAM(13689) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(13689))))  severity failure;
	assert RAM(13690) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(13690))))  severity failure;
	assert RAM(13691) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(13691))))  severity failure;
	assert RAM(13692) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(13692))))  severity failure;
	assert RAM(13693) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(13693))))  severity failure;
	assert RAM(13694) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(13694))))  severity failure;
	assert RAM(13695) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(13695))))  severity failure;
	assert RAM(13696) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(13696))))  severity failure;
	assert RAM(13697) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(13697))))  severity failure;
	assert RAM(13698) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(13698))))  severity failure;
	assert RAM(13699) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(13699))))  severity failure;
	assert RAM(13700) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(13700))))  severity failure;
	assert RAM(13701) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13701))))  severity failure;
	assert RAM(13702) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(13702))))  severity failure;
	assert RAM(13703) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(13703))))  severity failure;
	assert RAM(13704) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(13704))))  severity failure;
	assert RAM(13705) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(13705))))  severity failure;
	assert RAM(13706) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(13706))))  severity failure;
	assert RAM(13707) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(13707))))  severity failure;
	assert RAM(13708) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(13708))))  severity failure;
	assert RAM(13709) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(13709))))  severity failure;
	assert RAM(13710) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(13710))))  severity failure;
	assert RAM(13711) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(13711))))  severity failure;
	assert RAM(13712) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(13712))))  severity failure;
	assert RAM(13713) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(13713))))  severity failure;
	assert RAM(13714) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(13714))))  severity failure;
	assert RAM(13715) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(13715))))  severity failure;
	assert RAM(13716) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(13716))))  severity failure;
	assert RAM(13717) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(13717))))  severity failure;
	assert RAM(13718) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13718))))  severity failure;
	assert RAM(13719) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(13719))))  severity failure;
	assert RAM(13720) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(13720))))  severity failure;
	assert RAM(13721) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(13721))))  severity failure;
	assert RAM(13722) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(13722))))  severity failure;
	assert RAM(13723) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(13723))))  severity failure;
	assert RAM(13724) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(13724))))  severity failure;
	assert RAM(13725) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(13725))))  severity failure;
	assert RAM(13726) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(13726))))  severity failure;
	assert RAM(13727) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(13727))))  severity failure;
	assert RAM(13728) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(13728))))  severity failure;
	assert RAM(13729) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(13729))))  severity failure;
	assert RAM(13730) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(13730))))  severity failure;
	assert RAM(13731) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(13731))))  severity failure;
	assert RAM(13732) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(13732))))  severity failure;
	assert RAM(13733) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(13733))))  severity failure;
	assert RAM(13734) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(13734))))  severity failure;
	assert RAM(13735) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(13735))))  severity failure;
	assert RAM(13736) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(13736))))  severity failure;
	assert RAM(13737) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(13737))))  severity failure;
	assert RAM(13738) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(13738))))  severity failure;
	assert RAM(13739) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(13739))))  severity failure;
	assert RAM(13740) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(13740))))  severity failure;
	assert RAM(13741) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(13741))))  severity failure;
	assert RAM(13742) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(13742))))  severity failure;
	assert RAM(13743) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(13743))))  severity failure;
	assert RAM(13744) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(13744))))  severity failure;
	assert RAM(13745) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(13745))))  severity failure;
	assert RAM(13746) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(13746))))  severity failure;
	assert RAM(13747) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(13747))))  severity failure;
	assert RAM(13748) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(13748))))  severity failure;
	assert RAM(13749) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(13749))))  severity failure;
	assert RAM(13750) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(13750))))  severity failure;
	assert RAM(13751) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(13751))))  severity failure;
	assert RAM(13752) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(13752))))  severity failure;
	assert RAM(13753) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(13753))))  severity failure;
	assert RAM(13754) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(13754))))  severity failure;
	assert RAM(13755) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(13755))))  severity failure;
	assert RAM(13756) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(13756))))  severity failure;
	assert RAM(13757) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(13757))))  severity failure;
	assert RAM(13758) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(13758))))  severity failure;
	assert RAM(13759) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(13759))))  severity failure;
	assert RAM(13760) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(13760))))  severity failure;
	assert RAM(13761) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13761))))  severity failure;
	assert RAM(13762) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(13762))))  severity failure;
	assert RAM(13763) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(13763))))  severity failure;
	assert RAM(13764) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(13764))))  severity failure;
	assert RAM(13765) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(13765))))  severity failure;
	assert RAM(13766) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(13766))))  severity failure;
	assert RAM(13767) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(13767))))  severity failure;
	assert RAM(13768) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(13768))))  severity failure;
	assert RAM(13769) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(13769))))  severity failure;
	assert RAM(13770) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(13770))))  severity failure;
	assert RAM(13771) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(13771))))  severity failure;
	assert RAM(13772) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(13772))))  severity failure;
	assert RAM(13773) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(13773))))  severity failure;
	assert RAM(13774) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(13774))))  severity failure;
	assert RAM(13775) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(13775))))  severity failure;
	assert RAM(13776) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(13776))))  severity failure;
	assert RAM(13777) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(13777))))  severity failure;
	assert RAM(13778) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(13778))))  severity failure;
	assert RAM(13779) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(13779))))  severity failure;
	assert RAM(13780) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(13780))))  severity failure;
	assert RAM(13781) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(13781))))  severity failure;
	assert RAM(13782) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(13782))))  severity failure;
	assert RAM(13783) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(13783))))  severity failure;
	assert RAM(13784) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(13784))))  severity failure;
	assert RAM(13785) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(13785))))  severity failure;
	assert RAM(13786) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(13786))))  severity failure;
	assert RAM(13787) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(13787))))  severity failure;
	assert RAM(13788) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(13788))))  severity failure;
	assert RAM(13789) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(13789))))  severity failure;
	assert RAM(13790) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(13790))))  severity failure;
	assert RAM(13791) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(13791))))  severity failure;
	assert RAM(13792) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(13792))))  severity failure;
	assert RAM(13793) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(13793))))  severity failure;
	assert RAM(13794) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(13794))))  severity failure;
	assert RAM(13795) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(13795))))  severity failure;
	assert RAM(13796) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13796))))  severity failure;
	assert RAM(13797) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(13797))))  severity failure;
	assert RAM(13798) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(13798))))  severity failure;
	assert RAM(13799) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(13799))))  severity failure;
	assert RAM(13800) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(13800))))  severity failure;
	assert RAM(13801) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(13801))))  severity failure;
	assert RAM(13802) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(13802))))  severity failure;
	assert RAM(13803) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(13803))))  severity failure;
	assert RAM(13804) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(13804))))  severity failure;
	assert RAM(13805) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(13805))))  severity failure;
	assert RAM(13806) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(13806))))  severity failure;
	assert RAM(13807) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(13807))))  severity failure;
	assert RAM(13808) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(13808))))  severity failure;
	assert RAM(13809) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(13809))))  severity failure;
	assert RAM(13810) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(13810))))  severity failure;
	assert RAM(13811) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(13811))))  severity failure;
	assert RAM(13812) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(13812))))  severity failure;
	assert RAM(13813) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(13813))))  severity failure;
	assert RAM(13814) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(13814))))  severity failure;
	assert RAM(13815) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(13815))))  severity failure;
	assert RAM(13816) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(13816))))  severity failure;
	assert RAM(13817) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(13817))))  severity failure;
	assert RAM(13818) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(13818))))  severity failure;
	assert RAM(13819) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(13819))))  severity failure;
	assert RAM(13820) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(13820))))  severity failure;
	assert RAM(13821) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(13821))))  severity failure;
	assert RAM(13822) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(13822))))  severity failure;
	assert RAM(13823) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(13823))))  severity failure;
	assert RAM(13824) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(13824))))  severity failure;
	assert RAM(13825) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13825))))  severity failure;
	assert RAM(13826) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(13826))))  severity failure;
	assert RAM(13827) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(13827))))  severity failure;
	assert RAM(13828) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(13828))))  severity failure;
	assert RAM(13829) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(13829))))  severity failure;
	assert RAM(13830) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(13830))))  severity failure;
	assert RAM(13831) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(13831))))  severity failure;
	assert RAM(13832) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(13832))))  severity failure;
	assert RAM(13833) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(13833))))  severity failure;
	assert RAM(13834) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(13834))))  severity failure;
	assert RAM(13835) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(13835))))  severity failure;
	assert RAM(13836) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(13836))))  severity failure;
	assert RAM(13837) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(13837))))  severity failure;
	assert RAM(13838) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(13838))))  severity failure;
	assert RAM(13839) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(13839))))  severity failure;
	assert RAM(13840) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(13840))))  severity failure;
	assert RAM(13841) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(13841))))  severity failure;
	assert RAM(13842) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(13842))))  severity failure;
	assert RAM(13843) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(13843))))  severity failure;
	assert RAM(13844) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(13844))))  severity failure;
	assert RAM(13845) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(13845))))  severity failure;
	assert RAM(13846) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(13846))))  severity failure;
	assert RAM(13847) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(13847))))  severity failure;
	assert RAM(13848) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(13848))))  severity failure;
	assert RAM(13849) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13849))))  severity failure;
	assert RAM(13850) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(13850))))  severity failure;
	assert RAM(13851) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(13851))))  severity failure;
	assert RAM(13852) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13852))))  severity failure;
	assert RAM(13853) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(13853))))  severity failure;
	assert RAM(13854) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(13854))))  severity failure;
	assert RAM(13855) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(13855))))  severity failure;
	assert RAM(13856) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(13856))))  severity failure;
	assert RAM(13857) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(13857))))  severity failure;
	assert RAM(13858) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(13858))))  severity failure;
	assert RAM(13859) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(13859))))  severity failure;
	assert RAM(13860) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(13860))))  severity failure;
	assert RAM(13861) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(13861))))  severity failure;
	assert RAM(13862) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(13862))))  severity failure;
	assert RAM(13863) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(13863))))  severity failure;
	assert RAM(13864) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(13864))))  severity failure;
	assert RAM(13865) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(13865))))  severity failure;
	assert RAM(13866) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(13866))))  severity failure;
	assert RAM(13867) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(13867))))  severity failure;
	assert RAM(13868) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(13868))))  severity failure;
	assert RAM(13869) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(13869))))  severity failure;
	assert RAM(13870) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(13870))))  severity failure;
	assert RAM(13871) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(13871))))  severity failure;
	assert RAM(13872) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(13872))))  severity failure;
	assert RAM(13873) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(13873))))  severity failure;
	assert RAM(13874) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(13874))))  severity failure;
	assert RAM(13875) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(13875))))  severity failure;
	assert RAM(13876) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(13876))))  severity failure;
	assert RAM(13877) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(13877))))  severity failure;
	assert RAM(13878) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(13878))))  severity failure;
	assert RAM(13879) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(13879))))  severity failure;
	assert RAM(13880) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(13880))))  severity failure;
	assert RAM(13881) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(13881))))  severity failure;
	assert RAM(13882) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(13882))))  severity failure;
	assert RAM(13883) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(13883))))  severity failure;
	assert RAM(13884) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(13884))))  severity failure;
	assert RAM(13885) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(13885))))  severity failure;
	assert RAM(13886) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(13886))))  severity failure;
	assert RAM(13887) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(13887))))  severity failure;
	assert RAM(13888) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(13888))))  severity failure;
	assert RAM(13889) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(13889))))  severity failure;
	assert RAM(13890) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(13890))))  severity failure;
	assert RAM(13891) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(13891))))  severity failure;
	assert RAM(13892) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(13892))))  severity failure;
	assert RAM(13893) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(13893))))  severity failure;
	assert RAM(13894) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(13894))))  severity failure;
	assert RAM(13895) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(13895))))  severity failure;
	assert RAM(13896) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(13896))))  severity failure;
	assert RAM(13897) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(13897))))  severity failure;
	assert RAM(13898) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(13898))))  severity failure;
	assert RAM(13899) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(13899))))  severity failure;
	assert RAM(13900) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(13900))))  severity failure;
	assert RAM(13901) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(13901))))  severity failure;
	assert RAM(13902) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(13902))))  severity failure;
	assert RAM(13903) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(13903))))  severity failure;
	assert RAM(13904) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(13904))))  severity failure;
	assert RAM(13905) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(13905))))  severity failure;
	assert RAM(13906) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(13906))))  severity failure;
	assert RAM(13907) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(13907))))  severity failure;
	assert RAM(13908) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(13908))))  severity failure;
	assert RAM(13909) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(13909))))  severity failure;
	assert RAM(13910) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(13910))))  severity failure;
	assert RAM(13911) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(13911))))  severity failure;
	assert RAM(13912) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(13912))))  severity failure;
	assert RAM(13913) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(13913))))  severity failure;
	assert RAM(13914) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(13914))))  severity failure;
	assert RAM(13915) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(13915))))  severity failure;
	assert RAM(13916) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(13916))))  severity failure;
	assert RAM(13917) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(13917))))  severity failure;
	assert RAM(13918) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(13918))))  severity failure;
	assert RAM(13919) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(13919))))  severity failure;
	assert RAM(13920) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(13920))))  severity failure;
	assert RAM(13921) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(13921))))  severity failure;
	assert RAM(13922) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(13922))))  severity failure;
	assert RAM(13923) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(13923))))  severity failure;
	assert RAM(13924) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(13924))))  severity failure;
	assert RAM(13925) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(13925))))  severity failure;
	assert RAM(13926) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(13926))))  severity failure;
	assert RAM(13927) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(13927))))  severity failure;
	assert RAM(13928) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(13928))))  severity failure;
	assert RAM(13929) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(13929))))  severity failure;
	assert RAM(13930) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(13930))))  severity failure;
	assert RAM(13931) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(13931))))  severity failure;
	assert RAM(13932) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(13932))))  severity failure;
	assert RAM(13933) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(13933))))  severity failure;
	assert RAM(13934) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(13934))))  severity failure;
	assert RAM(13935) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(13935))))  severity failure;
	assert RAM(13936) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(13936))))  severity failure;
	assert RAM(13937) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(13937))))  severity failure;
	assert RAM(13938) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(13938))))  severity failure;
	assert RAM(13939) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(13939))))  severity failure;
	assert RAM(13940) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(13940))))  severity failure;
	assert RAM(13941) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(13941))))  severity failure;
	assert RAM(13942) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(13942))))  severity failure;
	assert RAM(13943) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(13943))))  severity failure;
	assert RAM(13944) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(13944))))  severity failure;
	assert RAM(13945) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(13945))))  severity failure;
	assert RAM(13946) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(13946))))  severity failure;
	assert RAM(13947) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(13947))))  severity failure;
	assert RAM(13948) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(13948))))  severity failure;
	assert RAM(13949) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(13949))))  severity failure;
	assert RAM(13950) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(13950))))  severity failure;
	assert RAM(13951) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(13951))))  severity failure;
	assert RAM(13952) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(13952))))  severity failure;
	assert RAM(13953) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(13953))))  severity failure;
	assert RAM(13954) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(13954))))  severity failure;
	assert RAM(13955) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(13955))))  severity failure;
	assert RAM(13956) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(13956))))  severity failure;
	assert RAM(13957) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(13957))))  severity failure;
	assert RAM(13958) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(13958))))  severity failure;
	assert RAM(13959) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(13959))))  severity failure;
	assert RAM(13960) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(13960))))  severity failure;
	assert RAM(13961) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(13961))))  severity failure;
	assert RAM(13962) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(13962))))  severity failure;
	assert RAM(13963) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(13963))))  severity failure;
	assert RAM(13964) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(13964))))  severity failure;
	assert RAM(13965) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(13965))))  severity failure;
	assert RAM(13966) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(13966))))  severity failure;
	assert RAM(13967) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(13967))))  severity failure;
	assert RAM(13968) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(13968))))  severity failure;
	assert RAM(13969) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(13969))))  severity failure;
	assert RAM(13970) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(13970))))  severity failure;
	assert RAM(13971) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(13971))))  severity failure;
	assert RAM(13972) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(13972))))  severity failure;
	assert RAM(13973) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(13973))))  severity failure;
	assert RAM(13974) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(13974))))  severity failure;
	assert RAM(13975) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(13975))))  severity failure;
	assert RAM(13976) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(13976))))  severity failure;
	assert RAM(13977) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(13977))))  severity failure;
	assert RAM(13978) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(13978))))  severity failure;
	assert RAM(13979) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(13979))))  severity failure;
	assert RAM(13980) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(13980))))  severity failure;
	assert RAM(13981) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(13981))))  severity failure;
	assert RAM(13982) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(13982))))  severity failure;
	assert RAM(13983) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(13983))))  severity failure;
	assert RAM(13984) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(13984))))  severity failure;
	assert RAM(13985) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(13985))))  severity failure;
	assert RAM(13986) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(13986))))  severity failure;
	assert RAM(13987) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(13987))))  severity failure;
	assert RAM(13988) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(13988))))  severity failure;
	assert RAM(13989) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(13989))))  severity failure;
	assert RAM(13990) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(13990))))  severity failure;
	assert RAM(13991) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(13991))))  severity failure;
	assert RAM(13992) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(13992))))  severity failure;
	assert RAM(13993) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(13993))))  severity failure;
	assert RAM(13994) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(13994))))  severity failure;
	assert RAM(13995) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(13995))))  severity failure;
	assert RAM(13996) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(13996))))  severity failure;
	assert RAM(13997) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(13997))))  severity failure;
	assert RAM(13998) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(13998))))  severity failure;
	assert RAM(13999) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(13999))))  severity failure;
	assert RAM(14000) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(14000))))  severity failure;
	assert RAM(14001) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(14001))))  severity failure;
	assert RAM(14002) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(14002))))  severity failure;
	assert RAM(14003) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(14003))))  severity failure;
	assert RAM(14004) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(14004))))  severity failure;
	assert RAM(14005) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(14005))))  severity failure;
	assert RAM(14006) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(14006))))  severity failure;
	assert RAM(14007) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(14007))))  severity failure;
	assert RAM(14008) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(14008))))  severity failure;
	assert RAM(14009) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(14009))))  severity failure;
	assert RAM(14010) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(14010))))  severity failure;
	assert RAM(14011) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(14011))))  severity failure;
	assert RAM(14012) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(14012))))  severity failure;
	assert RAM(14013) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(14013))))  severity failure;
	assert RAM(14014) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(14014))))  severity failure;
	assert RAM(14015) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(14015))))  severity failure;
	assert RAM(14016) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(14016))))  severity failure;
	assert RAM(14017) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(14017))))  severity failure;
	assert RAM(14018) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(14018))))  severity failure;
	assert RAM(14019) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(14019))))  severity failure;
	assert RAM(14020) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(14020))))  severity failure;
	assert RAM(14021) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(14021))))  severity failure;
	assert RAM(14022) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(14022))))  severity failure;
	assert RAM(14023) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(14023))))  severity failure;
	assert RAM(14024) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(14024))))  severity failure;
	assert RAM(14025) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(14025))))  severity failure;
	assert RAM(14026) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(14026))))  severity failure;
	assert RAM(14027) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(14027))))  severity failure;
	assert RAM(14028) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(14028))))  severity failure;
	assert RAM(14029) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(14029))))  severity failure;
	assert RAM(14030) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(14030))))  severity failure;
	assert RAM(14031) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(14031))))  severity failure;
	assert RAM(14032) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(14032))))  severity failure;
	assert RAM(14033) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(14033))))  severity failure;
	assert RAM(14034) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(14034))))  severity failure;
	assert RAM(14035) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(14035))))  severity failure;
	assert RAM(14036) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(14036))))  severity failure;
	assert RAM(14037) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(14037))))  severity failure;
	assert RAM(14038) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(14038))))  severity failure;
	assert RAM(14039) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(14039))))  severity failure;
	assert RAM(14040) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(14040))))  severity failure;
	assert RAM(14041) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(14041))))  severity failure;
	assert RAM(14042) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(14042))))  severity failure;
	assert RAM(14043) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(14043))))  severity failure;
	assert RAM(14044) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(14044))))  severity failure;
	assert RAM(14045) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(14045))))  severity failure;
	assert RAM(14046) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(14046))))  severity failure;
	assert RAM(14047) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(14047))))  severity failure;
	assert RAM(14048) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(14048))))  severity failure;
	assert RAM(14049) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(14049))))  severity failure;
	assert RAM(14050) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(14050))))  severity failure;
	assert RAM(14051) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(14051))))  severity failure;
	assert RAM(14052) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(14052))))  severity failure;
	assert RAM(14053) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(14053))))  severity failure;
	assert RAM(14054) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(14054))))  severity failure;
	assert RAM(14055) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(14055))))  severity failure;
	assert RAM(14056) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(14056))))  severity failure;
	assert RAM(14057) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(14057))))  severity failure;
	assert RAM(14058) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(14058))))  severity failure;
	assert RAM(14059) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(14059))))  severity failure;
	assert RAM(14060) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(14060))))  severity failure;
	assert RAM(14061) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(14061))))  severity failure;
	assert RAM(14062) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(14062))))  severity failure;
	assert RAM(14063) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(14063))))  severity failure;
	assert RAM(14064) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(14064))))  severity failure;
	assert RAM(14065) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(14065))))  severity failure;
	assert RAM(14066) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(14066))))  severity failure;
	assert RAM(14067) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(14067))))  severity failure;
	assert RAM(14068) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(14068))))  severity failure;
	assert RAM(14069) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(14069))))  severity failure;
	assert RAM(14070) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(14070))))  severity failure;
	assert RAM(14071) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(14071))))  severity failure;
	assert RAM(14072) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(14072))))  severity failure;
	assert RAM(14073) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(14073))))  severity failure;
	assert RAM(14074) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(14074))))  severity failure;
	assert RAM(14075) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(14075))))  severity failure;
	assert RAM(14076) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(14076))))  severity failure;
	assert RAM(14077) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(14077))))  severity failure;
	assert RAM(14078) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(14078))))  severity failure;
	assert RAM(14079) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(14079))))  severity failure;
	assert RAM(14080) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(14080))))  severity failure;
	assert RAM(14081) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(14081))))  severity failure;
	assert RAM(14082) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(14082))))  severity failure;
	assert RAM(14083) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(14083))))  severity failure;
	assert RAM(14084) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(14084))))  severity failure;
	assert RAM(14085) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(14085))))  severity failure;
	assert RAM(14086) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(14086))))  severity failure;
	assert RAM(14087) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(14087))))  severity failure;
	assert RAM(14088) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(14088))))  severity failure;
	assert RAM(14089) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(14089))))  severity failure;
	assert RAM(14090) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(14090))))  severity failure;
	assert RAM(14091) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(14091))))  severity failure;
	assert RAM(14092) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(14092))))  severity failure;
	assert RAM(14093) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(14093))))  severity failure;
	assert RAM(14094) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(14094))))  severity failure;
	assert RAM(14095) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(14095))))  severity failure;
	assert RAM(14096) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(14096))))  severity failure;
	assert RAM(14097) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(14097))))  severity failure;
	assert RAM(14098) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(14098))))  severity failure;
	assert RAM(14099) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(14099))))  severity failure;
	assert RAM(14100) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(14100))))  severity failure;
	assert RAM(14101) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(14101))))  severity failure;
	assert RAM(14102) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(14102))))  severity failure;
	assert RAM(14103) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(14103))))  severity failure;
	assert RAM(14104) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(14104))))  severity failure;
	assert RAM(14105) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(14105))))  severity failure;
	assert RAM(14106) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(14106))))  severity failure;
	assert RAM(14107) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(14107))))  severity failure;
	assert RAM(14108) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(14108))))  severity failure;
	assert RAM(14109) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(14109))))  severity failure;
	assert RAM(14110) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(14110))))  severity failure;
	assert RAM(14111) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(14111))))  severity failure;
	assert RAM(14112) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(14112))))  severity failure;
	assert RAM(14113) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(14113))))  severity failure;
	assert RAM(14114) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(14114))))  severity failure;
	assert RAM(14115) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(14115))))  severity failure;
	assert RAM(14116) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(14116))))  severity failure;
	assert RAM(14117) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(14117))))  severity failure;
	assert RAM(14118) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(14118))))  severity failure;
	assert RAM(14119) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(14119))))  severity failure;
	assert RAM(14120) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(14120))))  severity failure;
	assert RAM(14121) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(14121))))  severity failure;
	assert RAM(14122) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(14122))))  severity failure;
	assert RAM(14123) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(14123))))  severity failure;
	assert RAM(14124) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(14124))))  severity failure;
	assert RAM(14125) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(14125))))  severity failure;
	assert RAM(14126) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(14126))))  severity failure;
	assert RAM(14127) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(14127))))  severity failure;
	assert RAM(14128) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(14128))))  severity failure;
	assert RAM(14129) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(14129))))  severity failure;
	assert RAM(14130) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(14130))))  severity failure;
	assert RAM(14131) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(14131))))  severity failure;
	assert RAM(14132) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(14132))))  severity failure;
	assert RAM(14133) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(14133))))  severity failure;
	assert RAM(14134) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(14134))))  severity failure;
	assert RAM(14135) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(14135))))  severity failure;
	assert RAM(14136) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(14136))))  severity failure;
	assert RAM(14137) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(14137))))  severity failure;
	assert RAM(14138) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(14138))))  severity failure;
	assert RAM(14139) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(14139))))  severity failure;
	assert RAM(14140) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(14140))))  severity failure;
	assert RAM(14141) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(14141))))  severity failure;
	assert RAM(14142) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(14142))))  severity failure;
	assert RAM(14143) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(14143))))  severity failure;
	assert RAM(14144) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(14144))))  severity failure;
	assert RAM(14145) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(14145))))  severity failure;
	assert RAM(14146) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(14146))))  severity failure;
	assert RAM(14147) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(14147))))  severity failure;
	assert RAM(14148) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(14148))))  severity failure;
	assert RAM(14149) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(14149))))  severity failure;
	assert RAM(14150) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(14150))))  severity failure;
	assert RAM(14151) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(14151))))  severity failure;
	assert RAM(14152) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(14152))))  severity failure;
	assert RAM(14153) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(14153))))  severity failure;
	assert RAM(14154) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(14154))))  severity failure;
	assert RAM(14155) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(14155))))  severity failure;
	assert RAM(14156) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(14156))))  severity failure;
	assert RAM(14157) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(14157))))  severity failure;
	assert RAM(14158) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(14158))))  severity failure;
	assert RAM(14159) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(14159))))  severity failure;
	assert RAM(14160) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(14160))))  severity failure;
	assert RAM(14161) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(14161))))  severity failure;
	assert RAM(14162) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(14162))))  severity failure;
	assert RAM(14163) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(14163))))  severity failure;
	assert RAM(14164) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(14164))))  severity failure;
	assert RAM(14165) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(14165))))  severity failure;
	assert RAM(14166) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(14166))))  severity failure;
	assert RAM(14167) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(14167))))  severity failure;
	assert RAM(14168) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(14168))))  severity failure;
	assert RAM(14169) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(14169))))  severity failure;
	assert RAM(14170) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(14170))))  severity failure;
	assert RAM(14171) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(14171))))  severity failure;
	assert RAM(14172) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(14172))))  severity failure;
	assert RAM(14173) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(14173))))  severity failure;
	assert RAM(14174) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(14174))))  severity failure;
	assert RAM(14175) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(14175))))  severity failure;
	assert RAM(14176) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(14176))))  severity failure;
	assert RAM(14177) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(14177))))  severity failure;
	assert RAM(14178) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(14178))))  severity failure;
	assert RAM(14179) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(14179))))  severity failure;
	assert RAM(14180) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(14180))))  severity failure;
	assert RAM(14181) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(14181))))  severity failure;
	assert RAM(14182) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(14182))))  severity failure;
	assert RAM(14183) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(14183))))  severity failure;
	assert RAM(14184) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(14184))))  severity failure;
	assert RAM(14185) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(14185))))  severity failure;
	assert RAM(14186) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(14186))))  severity failure;
	assert RAM(14187) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(14187))))  severity failure;
	assert RAM(14188) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(14188))))  severity failure;
	assert RAM(14189) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(14189))))  severity failure;
	assert RAM(14190) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(14190))))  severity failure;
	assert RAM(14191) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(14191))))  severity failure;
	assert RAM(14192) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(14192))))  severity failure;
	assert RAM(14193) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(14193))))  severity failure;
	assert RAM(14194) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(14194))))  severity failure;
	assert RAM(14195) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(14195))))  severity failure;
	assert RAM(14196) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(14196))))  severity failure;
	assert RAM(14197) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(14197))))  severity failure;
	assert RAM(14198) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(14198))))  severity failure;
	assert RAM(14199) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(14199))))  severity failure;
	assert RAM(14200) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(14200))))  severity failure;
	assert RAM(14201) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(14201))))  severity failure;
	assert RAM(14202) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(14202))))  severity failure;
	assert RAM(14203) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(14203))))  severity failure;
	assert RAM(14204) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(14204))))  severity failure;
	assert RAM(14205) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(14205))))  severity failure;
	assert RAM(14206) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(14206))))  severity failure;
	assert RAM(14207) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(14207))))  severity failure;
	assert RAM(14208) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(14208))))  severity failure;
	assert RAM(14209) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(14209))))  severity failure;
	assert RAM(14210) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(14210))))  severity failure;
	assert RAM(14211) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(14211))))  severity failure;
	assert RAM(14212) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(14212))))  severity failure;
	assert RAM(14213) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(14213))))  severity failure;
	assert RAM(14214) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(14214))))  severity failure;
	assert RAM(14215) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(14215))))  severity failure;
	assert RAM(14216) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(14216))))  severity failure;
	assert RAM(14217) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(14217))))  severity failure;
	assert RAM(14218) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(14218))))  severity failure;
	assert RAM(14219) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(14219))))  severity failure;
	assert RAM(14220) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(14220))))  severity failure;
	assert RAM(14221) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(14221))))  severity failure;
	assert RAM(14222) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(14222))))  severity failure;
	assert RAM(14223) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(14223))))  severity failure;
	assert RAM(14224) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(14224))))  severity failure;
	assert RAM(14225) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(14225))))  severity failure;
	assert RAM(14226) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(14226))))  severity failure;
	assert RAM(14227) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(14227))))  severity failure;
	assert RAM(14228) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(14228))))  severity failure;
	assert RAM(14229) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(14229))))  severity failure;
	assert RAM(14230) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(14230))))  severity failure;
	assert RAM(14231) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(14231))))  severity failure;
	assert RAM(14232) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(14232))))  severity failure;
	assert RAM(14233) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(14233))))  severity failure;
	assert RAM(14234) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(14234))))  severity failure;
	assert RAM(14235) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(14235))))  severity failure;
	assert RAM(14236) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(14236))))  severity failure;
	assert RAM(14237) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(14237))))  severity failure;
	assert RAM(14238) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(14238))))  severity failure;
	assert RAM(14239) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(14239))))  severity failure;
	assert RAM(14240) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(14240))))  severity failure;
	assert RAM(14241) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(14241))))  severity failure;
	assert RAM(14242) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(14242))))  severity failure;
	assert RAM(14243) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(14243))))  severity failure;
	assert RAM(14244) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(14244))))  severity failure;
	assert RAM(14245) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(14245))))  severity failure;
	assert RAM(14246) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(14246))))  severity failure;
	assert RAM(14247) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(14247))))  severity failure;
	assert RAM(14248) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(14248))))  severity failure;
	assert RAM(14249) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(14249))))  severity failure;
	assert RAM(14250) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(14250))))  severity failure;
	assert RAM(14251) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(14251))))  severity failure;
	assert RAM(14252) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(14252))))  severity failure;
	assert RAM(14253) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(14253))))  severity failure;
	assert RAM(14254) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(14254))))  severity failure;
	assert RAM(14255) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(14255))))  severity failure;
	assert RAM(14256) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(14256))))  severity failure;
	assert RAM(14257) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(14257))))  severity failure;
	assert RAM(14258) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(14258))))  severity failure;
	assert RAM(14259) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(14259))))  severity failure;
	assert RAM(14260) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(14260))))  severity failure;
	assert RAM(14261) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(14261))))  severity failure;
	assert RAM(14262) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(14262))))  severity failure;
	assert RAM(14263) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(14263))))  severity failure;
	assert RAM(14264) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(14264))))  severity failure;
	assert RAM(14265) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(14265))))  severity failure;
	assert RAM(14266) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(14266))))  severity failure;
	assert RAM(14267) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(14267))))  severity failure;
	assert RAM(14268) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(14268))))  severity failure;
	assert RAM(14269) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(14269))))  severity failure;
	assert RAM(14270) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(14270))))  severity failure;
	assert RAM(14271) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(14271))))  severity failure;
	assert RAM(14272) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(14272))))  severity failure;
	assert RAM(14273) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(14273))))  severity failure;
	assert RAM(14274) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(14274))))  severity failure;
	assert RAM(14275) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(14275))))  severity failure;
	assert RAM(14276) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(14276))))  severity failure;
	assert RAM(14277) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(14277))))  severity failure;
	assert RAM(14278) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(14278))))  severity failure;
	assert RAM(14279) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(14279))))  severity failure;
	assert RAM(14280) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(14280))))  severity failure;
	assert RAM(14281) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(14281))))  severity failure;
	assert RAM(14282) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(14282))))  severity failure;
	assert RAM(14283) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(14283))))  severity failure;
	assert RAM(14284) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(14284))))  severity failure;
	assert RAM(14285) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(14285))))  severity failure;
	assert RAM(14286) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(14286))))  severity failure;
	assert RAM(14287) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(14287))))  severity failure;
	assert RAM(14288) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(14288))))  severity failure;
	assert RAM(14289) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(14289))))  severity failure;
	assert RAM(14290) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(14290))))  severity failure;
	assert RAM(14291) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(14291))))  severity failure;
	assert RAM(14292) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(14292))))  severity failure;
	assert RAM(14293) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(14293))))  severity failure;
	assert RAM(14294) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(14294))))  severity failure;
	assert RAM(14295) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(14295))))  severity failure;
	assert RAM(14296) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(14296))))  severity failure;
	assert RAM(14297) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(14297))))  severity failure;
	assert RAM(14298) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(14298))))  severity failure;
	assert RAM(14299) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(14299))))  severity failure;
	assert RAM(14300) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(14300))))  severity failure;
	assert RAM(14301) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(14301))))  severity failure;
	assert RAM(14302) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(14302))))  severity failure;
	assert RAM(14303) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(14303))))  severity failure;
	assert RAM(14304) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(14304))))  severity failure;
	assert RAM(14305) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(14305))))  severity failure;
	assert RAM(14306) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(14306))))  severity failure;
	assert RAM(14307) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(14307))))  severity failure;
	assert RAM(14308) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(14308))))  severity failure;
	assert RAM(14309) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(14309))))  severity failure;
	assert RAM(14310) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(14310))))  severity failure;
	assert RAM(14311) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(14311))))  severity failure;
	assert RAM(14312) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(14312))))  severity failure;
	assert RAM(14313) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(14313))))  severity failure;
	assert RAM(14314) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(14314))))  severity failure;
	assert RAM(14315) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(14315))))  severity failure;
	assert RAM(14316) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(14316))))  severity failure;
	assert RAM(14317) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(14317))))  severity failure;
	assert RAM(14318) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(14318))))  severity failure;
	assert RAM(14319) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(14319))))  severity failure;
	assert RAM(14320) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(14320))))  severity failure;
	assert RAM(14321) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(14321))))  severity failure;
	assert RAM(14322) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(14322))))  severity failure;
	assert RAM(14323) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(14323))))  severity failure;
	assert RAM(14324) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(14324))))  severity failure;
	assert RAM(14325) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(14325))))  severity failure;
	assert RAM(14326) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(14326))))  severity failure;
	assert RAM(14327) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(14327))))  severity failure;
	assert RAM(14328) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(14328))))  severity failure;
	assert RAM(14329) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(14329))))  severity failure;
	assert RAM(14330) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(14330))))  severity failure;
	assert RAM(14331) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(14331))))  severity failure;
	assert RAM(14332) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(14332))))  severity failure;
	assert RAM(14333) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(14333))))  severity failure;
	assert RAM(14334) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(14334))))  severity failure;
	assert RAM(14335) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(14335))))  severity failure;
	assert RAM(14336) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(14336))))  severity failure;
	assert RAM(14337) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(14337))))  severity failure;
	assert RAM(14338) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(14338))))  severity failure;
	assert RAM(14339) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(14339))))  severity failure;
	assert RAM(14340) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(14340))))  severity failure;
	assert RAM(14341) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(14341))))  severity failure;
	assert RAM(14342) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(14342))))  severity failure;
	assert RAM(14343) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(14343))))  severity failure;
	assert RAM(14344) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(14344))))  severity failure;
	assert RAM(14345) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(14345))))  severity failure;
	assert RAM(14346) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(14346))))  severity failure;
	assert RAM(14347) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(14347))))  severity failure;
	assert RAM(14348) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(14348))))  severity failure;
	assert RAM(14349) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(14349))))  severity failure;
	assert RAM(14350) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(14350))))  severity failure;
	assert RAM(14351) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(14351))))  severity failure;
	assert RAM(14352) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(14352))))  severity failure;
	assert RAM(14353) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(14353))))  severity failure;
	assert RAM(14354) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(14354))))  severity failure;
	assert RAM(14355) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(14355))))  severity failure;
	assert RAM(14356) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(14356))))  severity failure;
	assert RAM(14357) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(14357))))  severity failure;
	assert RAM(14358) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(14358))))  severity failure;
	assert RAM(14359) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(14359))))  severity failure;
	assert RAM(14360) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(14360))))  severity failure;
	assert RAM(14361) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(14361))))  severity failure;
	assert RAM(14362) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(14362))))  severity failure;
	assert RAM(14363) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(14363))))  severity failure;
	assert RAM(14364) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(14364))))  severity failure;
	assert RAM(14365) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(14365))))  severity failure;
	assert RAM(14366) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(14366))))  severity failure;
	assert RAM(14367) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(14367))))  severity failure;
	assert RAM(14368) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(14368))))  severity failure;
	assert RAM(14369) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(14369))))  severity failure;
	assert RAM(14370) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(14370))))  severity failure;
	assert RAM(14371) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(14371))))  severity failure;
	assert RAM(14372) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(14372))))  severity failure;
	assert RAM(14373) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(14373))))  severity failure;
	assert RAM(14374) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(14374))))  severity failure;
	assert RAM(14375) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(14375))))  severity failure;
	assert RAM(14376) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(14376))))  severity failure;
	assert RAM(14377) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(14377))))  severity failure;
	assert RAM(14378) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(14378))))  severity failure;
	assert RAM(14379) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(14379))))  severity failure;
	assert RAM(14380) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(14380))))  severity failure;
	assert RAM(14381) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(14381))))  severity failure;
	assert RAM(14382) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(14382))))  severity failure;
	assert RAM(14383) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(14383))))  severity failure;
	assert RAM(14384) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(14384))))  severity failure;
	assert RAM(14385) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(14385))))  severity failure;
	assert RAM(14386) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(14386))))  severity failure;
	assert RAM(14387) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(14387))))  severity failure;
	assert RAM(14388) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(14388))))  severity failure;
	assert RAM(14389) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(14389))))  severity failure;
	assert RAM(14390) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(14390))))  severity failure;
	assert RAM(14391) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(14391))))  severity failure;
	assert RAM(14392) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(14392))))  severity failure;
	assert RAM(14393) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(14393))))  severity failure;
	assert RAM(14394) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(14394))))  severity failure;
	assert RAM(14395) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(14395))))  severity failure;
	assert RAM(14396) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(14396))))  severity failure;
	assert RAM(14397) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(14397))))  severity failure;
	assert RAM(14398) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(14398))))  severity failure;
	assert RAM(14399) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(14399))))  severity failure;
	assert RAM(14400) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(14400))))  severity failure;
	assert RAM(14401) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(14401))))  severity failure;
	assert RAM(14402) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(14402))))  severity failure;
	assert RAM(14403) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(14403))))  severity failure;
	assert RAM(14404) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(14404))))  severity failure;
	assert RAM(14405) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(14405))))  severity failure;
	assert RAM(14406) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(14406))))  severity failure;
	assert RAM(14407) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(14407))))  severity failure;
	assert RAM(14408) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(14408))))  severity failure;
	assert RAM(14409) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(14409))))  severity failure;
	assert RAM(14410) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(14410))))  severity failure;
	assert RAM(14411) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(14411))))  severity failure;
	assert RAM(14412) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(14412))))  severity failure;
	assert RAM(14413) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(14413))))  severity failure;
	assert RAM(14414) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(14414))))  severity failure;
	assert RAM(14415) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(14415))))  severity failure;
	assert RAM(14416) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(14416))))  severity failure;
	assert RAM(14417) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(14417))))  severity failure;
	assert RAM(14418) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(14418))))  severity failure;
	assert RAM(14419) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(14419))))  severity failure;
	assert RAM(14420) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(14420))))  severity failure;
	assert RAM(14421) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(14421))))  severity failure;
	assert RAM(14422) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(14422))))  severity failure;
	assert RAM(14423) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(14423))))  severity failure;
	assert RAM(14424) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(14424))))  severity failure;
	assert RAM(14425) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(14425))))  severity failure;
	assert RAM(14426) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(14426))))  severity failure;
	assert RAM(14427) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(14427))))  severity failure;
	assert RAM(14428) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(14428))))  severity failure;
	assert RAM(14429) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(14429))))  severity failure;
	assert RAM(14430) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(14430))))  severity failure;
	assert RAM(14431) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(14431))))  severity failure;
	assert RAM(14432) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(14432))))  severity failure;
	assert RAM(14433) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(14433))))  severity failure;
	assert RAM(14434) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(14434))))  severity failure;
	assert RAM(14435) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(14435))))  severity failure;
	assert RAM(14436) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(14436))))  severity failure;
	assert RAM(14437) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(14437))))  severity failure;
	assert RAM(14438) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(14438))))  severity failure;
	assert RAM(14439) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(14439))))  severity failure;
	assert RAM(14440) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(14440))))  severity failure;
	assert RAM(14441) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(14441))))  severity failure;
	assert RAM(14442) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(14442))))  severity failure;
	assert RAM(14443) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(14443))))  severity failure;
	assert RAM(14444) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(14444))))  severity failure;
	assert RAM(14445) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(14445))))  severity failure;
	assert RAM(14446) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(14446))))  severity failure;
	assert RAM(14447) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(14447))))  severity failure;
	assert RAM(14448) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(14448))))  severity failure;
	assert RAM(14449) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(14449))))  severity failure;
	assert RAM(14450) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(14450))))  severity failure;
	assert RAM(14451) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(14451))))  severity failure;
	assert RAM(14452) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(14452))))  severity failure;
	assert RAM(14453) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(14453))))  severity failure;
	assert RAM(14454) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(14454))))  severity failure;
	assert RAM(14455) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(14455))))  severity failure;
	assert RAM(14456) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(14456))))  severity failure;
	assert RAM(14457) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(14457))))  severity failure;
	assert RAM(14458) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(14458))))  severity failure;
	assert RAM(14459) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(14459))))  severity failure;
	assert RAM(14460) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(14460))))  severity failure;
	assert RAM(14461) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(14461))))  severity failure;
	assert RAM(14462) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(14462))))  severity failure;
	assert RAM(14463) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(14463))))  severity failure;
	assert RAM(14464) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(14464))))  severity failure;
	assert RAM(14465) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(14465))))  severity failure;
	assert RAM(14466) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(14466))))  severity failure;
	assert RAM(14467) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(14467))))  severity failure;
	assert RAM(14468) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(14468))))  severity failure;
	assert RAM(14469) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(14469))))  severity failure;
	assert RAM(14470) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(14470))))  severity failure;
	assert RAM(14471) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(14471))))  severity failure;
	assert RAM(14472) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(14472))))  severity failure;
	assert RAM(14473) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(14473))))  severity failure;
	assert RAM(14474) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(14474))))  severity failure;
	assert RAM(14475) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(14475))))  severity failure;
	assert RAM(14476) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(14476))))  severity failure;
	assert RAM(14477) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(14477))))  severity failure;
	assert RAM(14478) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(14478))))  severity failure;
	assert RAM(14479) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(14479))))  severity failure;
	assert RAM(14480) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(14480))))  severity failure;
	assert RAM(14481) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(14481))))  severity failure;
	assert RAM(14482) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(14482))))  severity failure;
	assert RAM(14483) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(14483))))  severity failure;
	assert RAM(14484) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(14484))))  severity failure;
	assert RAM(14485) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(14485))))  severity failure;
	assert RAM(14486) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(14486))))  severity failure;
	assert RAM(14487) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(14487))))  severity failure;
	assert RAM(14488) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(14488))))  severity failure;
	assert RAM(14489) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(14489))))  severity failure;
	assert RAM(14490) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(14490))))  severity failure;
	assert RAM(14491) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(14491))))  severity failure;
	assert RAM(14492) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(14492))))  severity failure;
	assert RAM(14493) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(14493))))  severity failure;
	assert RAM(14494) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(14494))))  severity failure;
	assert RAM(14495) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(14495))))  severity failure;
	assert RAM(14496) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(14496))))  severity failure;
	assert RAM(14497) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(14497))))  severity failure;
	assert RAM(14498) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(14498))))  severity failure;
	assert RAM(14499) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(14499))))  severity failure;
	assert RAM(14500) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(14500))))  severity failure;
	assert RAM(14501) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(14501))))  severity failure;
	assert RAM(14502) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(14502))))  severity failure;
	assert RAM(14503) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(14503))))  severity failure;
	assert RAM(14504) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(14504))))  severity failure;
	assert RAM(14505) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(14505))))  severity failure;
	assert RAM(14506) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(14506))))  severity failure;
	assert RAM(14507) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(14507))))  severity failure;
	assert RAM(14508) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(14508))))  severity failure;
	assert RAM(14509) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(14509))))  severity failure;
	assert RAM(14510) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(14510))))  severity failure;
	assert RAM(14511) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(14511))))  severity failure;
	assert RAM(14512) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(14512))))  severity failure;
	assert RAM(14513) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(14513))))  severity failure;
	assert RAM(14514) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(14514))))  severity failure;
	assert RAM(14515) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(14515))))  severity failure;
	assert RAM(14516) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(14516))))  severity failure;
	assert RAM(14517) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(14517))))  severity failure;
	assert RAM(14518) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(14518))))  severity failure;
	assert RAM(14519) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(14519))))  severity failure;
	assert RAM(14520) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(14520))))  severity failure;
	assert RAM(14521) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(14521))))  severity failure;
	assert RAM(14522) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(14522))))  severity failure;
	assert RAM(14523) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(14523))))  severity failure;
	assert RAM(14524) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(14524))))  severity failure;
	assert RAM(14525) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(14525))))  severity failure;
	assert RAM(14526) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(14526))))  severity failure;
	assert RAM(14527) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(14527))))  severity failure;
	assert RAM(14528) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(14528))))  severity failure;
	assert RAM(14529) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(14529))))  severity failure;
	assert RAM(14530) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(14530))))  severity failure;
	assert RAM(14531) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(14531))))  severity failure;
	assert RAM(14532) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(14532))))  severity failure;
	assert RAM(14533) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(14533))))  severity failure;
	assert RAM(14534) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(14534))))  severity failure;
	assert RAM(14535) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(14535))))  severity failure;
	assert RAM(14536) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(14536))))  severity failure;
	assert RAM(14537) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(14537))))  severity failure;
	assert RAM(14538) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(14538))))  severity failure;
	assert RAM(14539) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(14539))))  severity failure;
	assert RAM(14540) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(14540))))  severity failure;
	assert RAM(14541) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(14541))))  severity failure;
	assert RAM(14542) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(14542))))  severity failure;
	assert RAM(14543) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(14543))))  severity failure;
	assert RAM(14544) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(14544))))  severity failure;
	assert RAM(14545) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(14545))))  severity failure;
	assert RAM(14546) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(14546))))  severity failure;
	assert RAM(14547) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(14547))))  severity failure;
	assert RAM(14548) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(14548))))  severity failure;
	assert RAM(14549) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(14549))))  severity failure;
	assert RAM(14550) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(14550))))  severity failure;
	assert RAM(14551) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(14551))))  severity failure;
	assert RAM(14552) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(14552))))  severity failure;
	assert RAM(14553) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(14553))))  severity failure;
	assert RAM(14554) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(14554))))  severity failure;
	assert RAM(14555) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(14555))))  severity failure;
	assert RAM(14556) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(14556))))  severity failure;
	assert RAM(14557) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(14557))))  severity failure;
	assert RAM(14558) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(14558))))  severity failure;
	assert RAM(14559) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(14559))))  severity failure;
	assert RAM(14560) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(14560))))  severity failure;
	assert RAM(14561) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(14561))))  severity failure;
	assert RAM(14562) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(14562))))  severity failure;
	assert RAM(14563) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(14563))))  severity failure;
	assert RAM(14564) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(14564))))  severity failure;
	assert RAM(14565) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(14565))))  severity failure;
	assert RAM(14566) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(14566))))  severity failure;
	assert RAM(14567) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(14567))))  severity failure;
	assert RAM(14568) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(14568))))  severity failure;
	assert RAM(14569) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(14569))))  severity failure;
	assert RAM(14570) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(14570))))  severity failure;
	assert RAM(14571) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(14571))))  severity failure;
	assert RAM(14572) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(14572))))  severity failure;
	assert RAM(14573) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(14573))))  severity failure;
	assert RAM(14574) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(14574))))  severity failure;
	assert RAM(14575) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(14575))))  severity failure;
	assert RAM(14576) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(14576))))  severity failure;
	assert RAM(14577) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(14577))))  severity failure;
	assert RAM(14578) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(14578))))  severity failure;
	assert RAM(14579) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(14579))))  severity failure;
	assert RAM(14580) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(14580))))  severity failure;
	assert RAM(14581) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(14581))))  severity failure;
	assert RAM(14582) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(14582))))  severity failure;
	assert RAM(14583) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(14583))))  severity failure;
	assert RAM(14584) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(14584))))  severity failure;
	assert RAM(14585) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(14585))))  severity failure;
	assert RAM(14586) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(14586))))  severity failure;
	assert RAM(14587) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(14587))))  severity failure;
	assert RAM(14588) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(14588))))  severity failure;
	assert RAM(14589) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(14589))))  severity failure;
	assert RAM(14590) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(14590))))  severity failure;
	assert RAM(14591) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(14591))))  severity failure;
	assert RAM(14592) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(14592))))  severity failure;
	assert RAM(14593) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(14593))))  severity failure;
	assert RAM(14594) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(14594))))  severity failure;
	assert RAM(14595) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(14595))))  severity failure;
	assert RAM(14596) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(14596))))  severity failure;
	assert RAM(14597) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(14597))))  severity failure;
	assert RAM(14598) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(14598))))  severity failure;
	assert RAM(14599) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(14599))))  severity failure;
	assert RAM(14600) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(14600))))  severity failure;
	assert RAM(14601) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(14601))))  severity failure;
	assert RAM(14602) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(14602))))  severity failure;
	assert RAM(14603) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(14603))))  severity failure;
	assert RAM(14604) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(14604))))  severity failure;
	assert RAM(14605) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(14605))))  severity failure;
	assert RAM(14606) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(14606))))  severity failure;
	assert RAM(14607) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(14607))))  severity failure;
	assert RAM(14608) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(14608))))  severity failure;
	assert RAM(14609) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(14609))))  severity failure;
	assert RAM(14610) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(14610))))  severity failure;
	assert RAM(14611) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(14611))))  severity failure;
	assert RAM(14612) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(14612))))  severity failure;
	assert RAM(14613) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(14613))))  severity failure;
	assert RAM(14614) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(14614))))  severity failure;
	assert RAM(14615) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(14615))))  severity failure;
	assert RAM(14616) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(14616))))  severity failure;
	assert RAM(14617) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(14617))))  severity failure;
	assert RAM(14618) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(14618))))  severity failure;
	assert RAM(14619) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(14619))))  severity failure;
	assert RAM(14620) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(14620))))  severity failure;
	assert RAM(14621) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(14621))))  severity failure;
	assert RAM(14622) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(14622))))  severity failure;
	assert RAM(14623) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(14623))))  severity failure;
	assert RAM(14624) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(14624))))  severity failure;
	assert RAM(14625) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(14625))))  severity failure;
	assert RAM(14626) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(14626))))  severity failure;
	assert RAM(14627) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(14627))))  severity failure;
	assert RAM(14628) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(14628))))  severity failure;
	assert RAM(14629) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(14629))))  severity failure;
	assert RAM(14630) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(14630))))  severity failure;
	assert RAM(14631) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(14631))))  severity failure;
	assert RAM(14632) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(14632))))  severity failure;
	assert RAM(14633) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(14633))))  severity failure;
	assert RAM(14634) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(14634))))  severity failure;
	assert RAM(14635) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(14635))))  severity failure;
	assert RAM(14636) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(14636))))  severity failure;
	assert RAM(14637) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(14637))))  severity failure;
	assert RAM(14638) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(14638))))  severity failure;
	assert RAM(14639) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(14639))))  severity failure;
	assert RAM(14640) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(14640))))  severity failure;
	assert RAM(14641) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(14641))))  severity failure;
	assert RAM(14642) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(14642))))  severity failure;
	assert RAM(14643) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(14643))))  severity failure;
	assert RAM(14644) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(14644))))  severity failure;
	assert RAM(14645) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(14645))))  severity failure;
	assert RAM(14646) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(14646))))  severity failure;
	assert RAM(14647) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(14647))))  severity failure;
	assert RAM(14648) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(14648))))  severity failure;
	assert RAM(14649) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(14649))))  severity failure;
	assert RAM(14650) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(14650))))  severity failure;
	assert RAM(14651) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(14651))))  severity failure;
	assert RAM(14652) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(14652))))  severity failure;
	assert RAM(14653) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(14653))))  severity failure;
	assert RAM(14654) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(14654))))  severity failure;
	assert RAM(14655) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(14655))))  severity failure;
	assert RAM(14656) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(14656))))  severity failure;
	assert RAM(14657) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(14657))))  severity failure;
	assert RAM(14658) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(14658))))  severity failure;
	assert RAM(14659) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(14659))))  severity failure;
	assert RAM(14660) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(14660))))  severity failure;
	assert RAM(14661) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(14661))))  severity failure;
	assert RAM(14662) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(14662))))  severity failure;
	assert RAM(14663) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(14663))))  severity failure;
	assert RAM(14664) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(14664))))  severity failure;
	assert RAM(14665) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(14665))))  severity failure;
	assert RAM(14666) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(14666))))  severity failure;
	assert RAM(14667) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(14667))))  severity failure;
	assert RAM(14668) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(14668))))  severity failure;
	assert RAM(14669) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(14669))))  severity failure;
	assert RAM(14670) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(14670))))  severity failure;
	assert RAM(14671) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(14671))))  severity failure;
	assert RAM(14672) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(14672))))  severity failure;
	assert RAM(14673) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(14673))))  severity failure;
	assert RAM(14674) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(14674))))  severity failure;
	assert RAM(14675) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(14675))))  severity failure;
	assert RAM(14676) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(14676))))  severity failure;
	assert RAM(14677) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(14677))))  severity failure;
	assert RAM(14678) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(14678))))  severity failure;
	assert RAM(14679) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(14679))))  severity failure;
	assert RAM(14680) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(14680))))  severity failure;
	assert RAM(14681) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(14681))))  severity failure;
	assert RAM(14682) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(14682))))  severity failure;
	assert RAM(14683) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(14683))))  severity failure;
	assert RAM(14684) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(14684))))  severity failure;
	assert RAM(14685) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(14685))))  severity failure;
	assert RAM(14686) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(14686))))  severity failure;
	assert RAM(14687) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(14687))))  severity failure;
	assert RAM(14688) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(14688))))  severity failure;
	assert RAM(14689) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(14689))))  severity failure;
	assert RAM(14690) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(14690))))  severity failure;
	assert RAM(14691) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(14691))))  severity failure;
	assert RAM(14692) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(14692))))  severity failure;
	assert RAM(14693) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(14693))))  severity failure;
	assert RAM(14694) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(14694))))  severity failure;
	assert RAM(14695) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(14695))))  severity failure;
	assert RAM(14696) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(14696))))  severity failure;
	assert RAM(14697) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(14697))))  severity failure;
	assert RAM(14698) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(14698))))  severity failure;
	assert RAM(14699) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(14699))))  severity failure;
	assert RAM(14700) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(14700))))  severity failure;
	assert RAM(14701) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(14701))))  severity failure;
	assert RAM(14702) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(14702))))  severity failure;
	assert RAM(14703) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(14703))))  severity failure;
	assert RAM(14704) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(14704))))  severity failure;
	assert RAM(14705) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(14705))))  severity failure;
	assert RAM(14706) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(14706))))  severity failure;
	assert RAM(14707) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(14707))))  severity failure;
	assert RAM(14708) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(14708))))  severity failure;
	assert RAM(14709) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(14709))))  severity failure;
	assert RAM(14710) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(14710))))  severity failure;
	assert RAM(14711) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(14711))))  severity failure;
	assert RAM(14712) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(14712))))  severity failure;
	assert RAM(14713) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(14713))))  severity failure;
	assert RAM(14714) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(14714))))  severity failure;
	assert RAM(14715) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(14715))))  severity failure;
	assert RAM(14716) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(14716))))  severity failure;
	assert RAM(14717) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(14717))))  severity failure;
	assert RAM(14718) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(14718))))  severity failure;
	assert RAM(14719) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(14719))))  severity failure;
	assert RAM(14720) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(14720))))  severity failure;
	assert RAM(14721) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(14721))))  severity failure;
	assert RAM(14722) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(14722))))  severity failure;
	assert RAM(14723) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(14723))))  severity failure;
	assert RAM(14724) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(14724))))  severity failure;
	assert RAM(14725) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(14725))))  severity failure;
	assert RAM(14726) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(14726))))  severity failure;
	assert RAM(14727) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(14727))))  severity failure;
	assert RAM(14728) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(14728))))  severity failure;
	assert RAM(14729) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(14729))))  severity failure;
	assert RAM(14730) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(14730))))  severity failure;
	assert RAM(14731) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(14731))))  severity failure;
	assert RAM(14732) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(14732))))  severity failure;
	assert RAM(14733) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(14733))))  severity failure;
	assert RAM(14734) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(14734))))  severity failure;
	assert RAM(14735) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(14735))))  severity failure;
	assert RAM(14736) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(14736))))  severity failure;
	assert RAM(14737) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(14737))))  severity failure;
	assert RAM(14738) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(14738))))  severity failure;
	assert RAM(14739) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(14739))))  severity failure;
	assert RAM(14740) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(14740))))  severity failure;
	assert RAM(14741) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(14741))))  severity failure;
	assert RAM(14742) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(14742))))  severity failure;
	assert RAM(14743) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(14743))))  severity failure;
	assert RAM(14744) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(14744))))  severity failure;
	assert RAM(14745) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(14745))))  severity failure;
	assert RAM(14746) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(14746))))  severity failure;
	assert RAM(14747) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(14747))))  severity failure;
	assert RAM(14748) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(14748))))  severity failure;
	assert RAM(14749) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(14749))))  severity failure;
	assert RAM(14750) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(14750))))  severity failure;
	assert RAM(14751) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(14751))))  severity failure;
	assert RAM(14752) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(14752))))  severity failure;
	assert RAM(14753) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(14753))))  severity failure;
	assert RAM(14754) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(14754))))  severity failure;
	assert RAM(14755) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(14755))))  severity failure;
	assert RAM(14756) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(14756))))  severity failure;
	assert RAM(14757) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(14757))))  severity failure;
	assert RAM(14758) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(14758))))  severity failure;
	assert RAM(14759) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(14759))))  severity failure;
	assert RAM(14760) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(14760))))  severity failure;
	assert RAM(14761) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(14761))))  severity failure;
	assert RAM(14762) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(14762))))  severity failure;
	assert RAM(14763) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(14763))))  severity failure;
	assert RAM(14764) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(14764))))  severity failure;
	assert RAM(14765) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(14765))))  severity failure;
	assert RAM(14766) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(14766))))  severity failure;
	assert RAM(14767) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(14767))))  severity failure;
	assert RAM(14768) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(14768))))  severity failure;
	assert RAM(14769) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(14769))))  severity failure;
	assert RAM(14770) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(14770))))  severity failure;
	assert RAM(14771) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(14771))))  severity failure;
	assert RAM(14772) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(14772))))  severity failure;
	assert RAM(14773) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(14773))))  severity failure;
	assert RAM(14774) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(14774))))  severity failure;
	assert RAM(14775) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(14775))))  severity failure;
	assert RAM(14776) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(14776))))  severity failure;
	assert RAM(14777) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(14777))))  severity failure;
	assert RAM(14778) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(14778))))  severity failure;
	assert RAM(14779) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(14779))))  severity failure;
	assert RAM(14780) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(14780))))  severity failure;
	assert RAM(14781) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(14781))))  severity failure;
	assert RAM(14782) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(14782))))  severity failure;
	assert RAM(14783) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(14783))))  severity failure;
	assert RAM(14784) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(14784))))  severity failure;
	assert RAM(14785) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(14785))))  severity failure;
	assert RAM(14786) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(14786))))  severity failure;
	assert RAM(14787) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(14787))))  severity failure;
	assert RAM(14788) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(14788))))  severity failure;
	assert RAM(14789) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(14789))))  severity failure;
	assert RAM(14790) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(14790))))  severity failure;
	assert RAM(14791) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(14791))))  severity failure;
	assert RAM(14792) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(14792))))  severity failure;
	assert RAM(14793) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(14793))))  severity failure;
	assert RAM(14794) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(14794))))  severity failure;
	assert RAM(14795) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(14795))))  severity failure;
	assert RAM(14796) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(14796))))  severity failure;
	assert RAM(14797) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(14797))))  severity failure;
	assert RAM(14798) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(14798))))  severity failure;
	assert RAM(14799) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(14799))))  severity failure;
	assert RAM(14800) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(14800))))  severity failure;
	assert RAM(14801) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(14801))))  severity failure;
	assert RAM(14802) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(14802))))  severity failure;
	assert RAM(14803) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(14803))))  severity failure;
	assert RAM(14804) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(14804))))  severity failure;
	assert RAM(14805) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(14805))))  severity failure;
	assert RAM(14806) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(14806))))  severity failure;
	assert RAM(14807) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(14807))))  severity failure;
	assert RAM(14808) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(14808))))  severity failure;
	assert RAM(14809) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(14809))))  severity failure;
	assert RAM(14810) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(14810))))  severity failure;
	assert RAM(14811) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(14811))))  severity failure;
	assert RAM(14812) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(14812))))  severity failure;
	assert RAM(14813) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(14813))))  severity failure;
	assert RAM(14814) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(14814))))  severity failure;
	assert RAM(14815) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(14815))))  severity failure;
	assert RAM(14816) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(14816))))  severity failure;
	assert RAM(14817) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(14817))))  severity failure;
	assert RAM(14818) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(14818))))  severity failure;
	assert RAM(14819) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(14819))))  severity failure;
	assert RAM(14820) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(14820))))  severity failure;
	assert RAM(14821) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(14821))))  severity failure;
	assert RAM(14822) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(14822))))  severity failure;
	assert RAM(14823) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(14823))))  severity failure;
	assert RAM(14824) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(14824))))  severity failure;
	assert RAM(14825) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(14825))))  severity failure;
	assert RAM(14826) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(14826))))  severity failure;
	assert RAM(14827) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(14827))))  severity failure;
	assert RAM(14828) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(14828))))  severity failure;
	assert RAM(14829) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(14829))))  severity failure;
	assert RAM(14830) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(14830))))  severity failure;
	assert RAM(14831) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(14831))))  severity failure;
	assert RAM(14832) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(14832))))  severity failure;
	assert RAM(14833) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(14833))))  severity failure;
	assert RAM(14834) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(14834))))  severity failure;
	assert RAM(14835) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(14835))))  severity failure;
	assert RAM(14836) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(14836))))  severity failure;
	assert RAM(14837) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(14837))))  severity failure;
	assert RAM(14838) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(14838))))  severity failure;
	assert RAM(14839) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(14839))))  severity failure;
	assert RAM(14840) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(14840))))  severity failure;
	assert RAM(14841) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(14841))))  severity failure;
	assert RAM(14842) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(14842))))  severity failure;
	assert RAM(14843) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(14843))))  severity failure;
	assert RAM(14844) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(14844))))  severity failure;
	assert RAM(14845) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(14845))))  severity failure;
	assert RAM(14846) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(14846))))  severity failure;
	assert RAM(14847) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(14847))))  severity failure;
	assert RAM(14848) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(14848))))  severity failure;
	assert RAM(14849) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(14849))))  severity failure;
	assert RAM(14850) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(14850))))  severity failure;
	assert RAM(14851) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(14851))))  severity failure;
	assert RAM(14852) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(14852))))  severity failure;
	assert RAM(14853) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(14853))))  severity failure;
	assert RAM(14854) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(14854))))  severity failure;
	assert RAM(14855) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(14855))))  severity failure;
	assert RAM(14856) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(14856))))  severity failure;
	assert RAM(14857) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(14857))))  severity failure;
	assert RAM(14858) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(14858))))  severity failure;
	assert RAM(14859) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(14859))))  severity failure;
	assert RAM(14860) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(14860))))  severity failure;
	assert RAM(14861) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(14861))))  severity failure;
	assert RAM(14862) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(14862))))  severity failure;
	assert RAM(14863) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(14863))))  severity failure;
	assert RAM(14864) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(14864))))  severity failure;
	assert RAM(14865) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(14865))))  severity failure;
	assert RAM(14866) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(14866))))  severity failure;
	assert RAM(14867) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(14867))))  severity failure;
	assert RAM(14868) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(14868))))  severity failure;
	assert RAM(14869) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(14869))))  severity failure;
	assert RAM(14870) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(14870))))  severity failure;
	assert RAM(14871) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(14871))))  severity failure;
	assert RAM(14872) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(14872))))  severity failure;
	assert RAM(14873) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(14873))))  severity failure;
	assert RAM(14874) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(14874))))  severity failure;
	assert RAM(14875) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(14875))))  severity failure;
	assert RAM(14876) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(14876))))  severity failure;
	assert RAM(14877) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(14877))))  severity failure;
	assert RAM(14878) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(14878))))  severity failure;
	assert RAM(14879) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(14879))))  severity failure;
	assert RAM(14880) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(14880))))  severity failure;
	assert RAM(14881) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(14881))))  severity failure;
	assert RAM(14882) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(14882))))  severity failure;
	assert RAM(14883) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(14883))))  severity failure;
	assert RAM(14884) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(14884))))  severity failure;
	assert RAM(14885) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(14885))))  severity failure;
	assert RAM(14886) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(14886))))  severity failure;
	assert RAM(14887) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(14887))))  severity failure;
	assert RAM(14888) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(14888))))  severity failure;
	assert RAM(14889) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(14889))))  severity failure;
	assert RAM(14890) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(14890))))  severity failure;
	assert RAM(14891) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(14891))))  severity failure;
	assert RAM(14892) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(14892))))  severity failure;
	assert RAM(14893) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(14893))))  severity failure;
	assert RAM(14894) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(14894))))  severity failure;
	assert RAM(14895) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(14895))))  severity failure;
	assert RAM(14896) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(14896))))  severity failure;
	assert RAM(14897) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(14897))))  severity failure;
	assert RAM(14898) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(14898))))  severity failure;
	assert RAM(14899) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(14899))))  severity failure;
	assert RAM(14900) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(14900))))  severity failure;
	assert RAM(14901) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(14901))))  severity failure;
	assert RAM(14902) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(14902))))  severity failure;
	assert RAM(14903) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(14903))))  severity failure;
	assert RAM(14904) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(14904))))  severity failure;
	assert RAM(14905) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(14905))))  severity failure;
	assert RAM(14906) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(14906))))  severity failure;
	assert RAM(14907) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(14907))))  severity failure;
	assert RAM(14908) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(14908))))  severity failure;
	assert RAM(14909) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(14909))))  severity failure;
	assert RAM(14910) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(14910))))  severity failure;
	assert RAM(14911) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(14911))))  severity failure;
	assert RAM(14912) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(14912))))  severity failure;
	assert RAM(14913) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(14913))))  severity failure;
	assert RAM(14914) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(14914))))  severity failure;
	assert RAM(14915) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(14915))))  severity failure;
	assert RAM(14916) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(14916))))  severity failure;
	assert RAM(14917) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(14917))))  severity failure;
	assert RAM(14918) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(14918))))  severity failure;
	assert RAM(14919) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(14919))))  severity failure;
	assert RAM(14920) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(14920))))  severity failure;
	assert RAM(14921) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(14921))))  severity failure;
	assert RAM(14922) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(14922))))  severity failure;
	assert RAM(14923) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(14923))))  severity failure;
	assert RAM(14924) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(14924))))  severity failure;
	assert RAM(14925) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(14925))))  severity failure;
	assert RAM(14926) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(14926))))  severity failure;
	assert RAM(14927) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(14927))))  severity failure;
	assert RAM(14928) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(14928))))  severity failure;
	assert RAM(14929) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(14929))))  severity failure;
	assert RAM(14930) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(14930))))  severity failure;
	assert RAM(14931) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(14931))))  severity failure;
	assert RAM(14932) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(14932))))  severity failure;
	assert RAM(14933) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(14933))))  severity failure;
	assert RAM(14934) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(14934))))  severity failure;
	assert RAM(14935) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(14935))))  severity failure;
	assert RAM(14936) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(14936))))  severity failure;
	assert RAM(14937) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(14937))))  severity failure;
	assert RAM(14938) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(14938))))  severity failure;
	assert RAM(14939) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(14939))))  severity failure;
	assert RAM(14940) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(14940))))  severity failure;
	assert RAM(14941) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(14941))))  severity failure;
	assert RAM(14942) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(14942))))  severity failure;
	assert RAM(14943) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(14943))))  severity failure;
	assert RAM(14944) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(14944))))  severity failure;
	assert RAM(14945) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(14945))))  severity failure;
	assert RAM(14946) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(14946))))  severity failure;
	assert RAM(14947) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(14947))))  severity failure;
	assert RAM(14948) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(14948))))  severity failure;
	assert RAM(14949) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(14949))))  severity failure;
	assert RAM(14950) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(14950))))  severity failure;
	assert RAM(14951) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(14951))))  severity failure;
	assert RAM(14952) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(14952))))  severity failure;
	assert RAM(14953) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(14953))))  severity failure;
	assert RAM(14954) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(14954))))  severity failure;
	assert RAM(14955) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(14955))))  severity failure;
	assert RAM(14956) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(14956))))  severity failure;
	assert RAM(14957) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(14957))))  severity failure;
	assert RAM(14958) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(14958))))  severity failure;
	assert RAM(14959) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(14959))))  severity failure;
	assert RAM(14960) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(14960))))  severity failure;
	assert RAM(14961) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(14961))))  severity failure;
	assert RAM(14962) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(14962))))  severity failure;
	assert RAM(14963) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(14963))))  severity failure;
	assert RAM(14964) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(14964))))  severity failure;
	assert RAM(14965) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(14965))))  severity failure;
	assert RAM(14966) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(14966))))  severity failure;
	assert RAM(14967) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(14967))))  severity failure;
	assert RAM(14968) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(14968))))  severity failure;
	assert RAM(14969) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(14969))))  severity failure;
	assert RAM(14970) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(14970))))  severity failure;
	assert RAM(14971) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(14971))))  severity failure;
	assert RAM(14972) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(14972))))  severity failure;
	assert RAM(14973) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(14973))))  severity failure;
	assert RAM(14974) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(14974))))  severity failure;
	assert RAM(14975) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(14975))))  severity failure;
	assert RAM(14976) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(14976))))  severity failure;
	assert RAM(14977) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(14977))))  severity failure;
	assert RAM(14978) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(14978))))  severity failure;
	assert RAM(14979) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(14979))))  severity failure;
	assert RAM(14980) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(14980))))  severity failure;
	assert RAM(14981) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(14981))))  severity failure;
	assert RAM(14982) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(14982))))  severity failure;
	assert RAM(14983) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(14983))))  severity failure;
	assert RAM(14984) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(14984))))  severity failure;
	assert RAM(14985) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(14985))))  severity failure;
	assert RAM(14986) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(14986))))  severity failure;
	assert RAM(14987) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(14987))))  severity failure;
	assert RAM(14988) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(14988))))  severity failure;
	assert RAM(14989) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(14989))))  severity failure;
	assert RAM(14990) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(14990))))  severity failure;
	assert RAM(14991) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(14991))))  severity failure;
	assert RAM(14992) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(14992))))  severity failure;
	assert RAM(14993) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(14993))))  severity failure;
	assert RAM(14994) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(14994))))  severity failure;
	assert RAM(14995) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(14995))))  severity failure;
	assert RAM(14996) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(14996))))  severity failure;
	assert RAM(14997) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(14997))))  severity failure;
	assert RAM(14998) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(14998))))  severity failure;
	assert RAM(14999) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(14999))))  severity failure;
	assert RAM(15000) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(15000))))  severity failure;
	assert RAM(15001) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(15001))))  severity failure;
	assert RAM(15002) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(15002))))  severity failure;
	assert RAM(15003) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(15003))))  severity failure;
	assert RAM(15004) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(15004))))  severity failure;
	assert RAM(15005) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(15005))))  severity failure;
	assert RAM(15006) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(15006))))  severity failure;
	assert RAM(15007) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(15007))))  severity failure;
	assert RAM(15008) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(15008))))  severity failure;
	assert RAM(15009) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(15009))))  severity failure;
	assert RAM(15010) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(15010))))  severity failure;
	assert RAM(15011) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(15011))))  severity failure;
	assert RAM(15012) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(15012))))  severity failure;
	assert RAM(15013) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(15013))))  severity failure;
	assert RAM(15014) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(15014))))  severity failure;
	assert RAM(15015) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(15015))))  severity failure;
	assert RAM(15016) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(15016))))  severity failure;
	assert RAM(15017) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(15017))))  severity failure;
	assert RAM(15018) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(15018))))  severity failure;
	assert RAM(15019) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(15019))))  severity failure;
	assert RAM(15020) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(15020))))  severity failure;
	assert RAM(15021) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(15021))))  severity failure;
	assert RAM(15022) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(15022))))  severity failure;
	assert RAM(15023) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(15023))))  severity failure;
	assert RAM(15024) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(15024))))  severity failure;
	assert RAM(15025) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(15025))))  severity failure;
	assert RAM(15026) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(15026))))  severity failure;
	assert RAM(15027) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(15027))))  severity failure;
	assert RAM(15028) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(15028))))  severity failure;
	assert RAM(15029) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(15029))))  severity failure;
	assert RAM(15030) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(15030))))  severity failure;
	assert RAM(15031) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(15031))))  severity failure;
	assert RAM(15032) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(15032))))  severity failure;
	assert RAM(15033) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(15033))))  severity failure;
	assert RAM(15034) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(15034))))  severity failure;
	assert RAM(15035) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(15035))))  severity failure;
	assert RAM(15036) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(15036))))  severity failure;
	assert RAM(15037) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(15037))))  severity failure;
	assert RAM(15038) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(15038))))  severity failure;
	assert RAM(15039) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(15039))))  severity failure;
	assert RAM(15040) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(15040))))  severity failure;
	assert RAM(15041) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(15041))))  severity failure;
	assert RAM(15042) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(15042))))  severity failure;
	assert RAM(15043) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(15043))))  severity failure;
	assert RAM(15044) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(15044))))  severity failure;
	assert RAM(15045) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(15045))))  severity failure;
	assert RAM(15046) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(15046))))  severity failure;
	assert RAM(15047) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(15047))))  severity failure;
	assert RAM(15048) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(15048))))  severity failure;
	assert RAM(15049) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(15049))))  severity failure;
	assert RAM(15050) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(15050))))  severity failure;
	assert RAM(15051) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15051))))  severity failure;
	assert RAM(15052) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(15052))))  severity failure;
	assert RAM(15053) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(15053))))  severity failure;
	assert RAM(15054) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(15054))))  severity failure;
	assert RAM(15055) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(15055))))  severity failure;
	assert RAM(15056) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(15056))))  severity failure;
	assert RAM(15057) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(15057))))  severity failure;
	assert RAM(15058) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(15058))))  severity failure;
	assert RAM(15059) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(15059))))  severity failure;
	assert RAM(15060) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(15060))))  severity failure;
	assert RAM(15061) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(15061))))  severity failure;
	assert RAM(15062) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(15062))))  severity failure;
	assert RAM(15063) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(15063))))  severity failure;
	assert RAM(15064) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(15064))))  severity failure;
	assert RAM(15065) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(15065))))  severity failure;
	assert RAM(15066) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(15066))))  severity failure;
	assert RAM(15067) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(15067))))  severity failure;
	assert RAM(15068) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(15068))))  severity failure;
	assert RAM(15069) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(15069))))  severity failure;
	assert RAM(15070) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(15070))))  severity failure;
	assert RAM(15071) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(15071))))  severity failure;
	assert RAM(15072) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(15072))))  severity failure;
	assert RAM(15073) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(15073))))  severity failure;
	assert RAM(15074) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(15074))))  severity failure;
	assert RAM(15075) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(15075))))  severity failure;
	assert RAM(15076) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(15076))))  severity failure;
	assert RAM(15077) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(15077))))  severity failure;
	assert RAM(15078) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(15078))))  severity failure;
	assert RAM(15079) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(15079))))  severity failure;
	assert RAM(15080) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(15080))))  severity failure;
	assert RAM(15081) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15081))))  severity failure;
	assert RAM(15082) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(15082))))  severity failure;
	assert RAM(15083) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(15083))))  severity failure;
	assert RAM(15084) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(15084))))  severity failure;
	assert RAM(15085) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(15085))))  severity failure;
	assert RAM(15086) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(15086))))  severity failure;
	assert RAM(15087) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(15087))))  severity failure;
	assert RAM(15088) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(15088))))  severity failure;
	assert RAM(15089) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(15089))))  severity failure;
	assert RAM(15090) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(15090))))  severity failure;
	assert RAM(15091) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(15091))))  severity failure;
	assert RAM(15092) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(15092))))  severity failure;
	assert RAM(15093) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(15093))))  severity failure;
	assert RAM(15094) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(15094))))  severity failure;
	assert RAM(15095) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(15095))))  severity failure;
	assert RAM(15096) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(15096))))  severity failure;
	assert RAM(15097) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(15097))))  severity failure;
	assert RAM(15098) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(15098))))  severity failure;
	assert RAM(15099) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(15099))))  severity failure;
	assert RAM(15100) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(15100))))  severity failure;
	assert RAM(15101) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(15101))))  severity failure;
	assert RAM(15102) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(15102))))  severity failure;
	assert RAM(15103) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(15103))))  severity failure;
	assert RAM(15104) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(15104))))  severity failure;
	assert RAM(15105) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(15105))))  severity failure;
	assert RAM(15106) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(15106))))  severity failure;
	assert RAM(15107) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(15107))))  severity failure;
	assert RAM(15108) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(15108))))  severity failure;
	assert RAM(15109) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(15109))))  severity failure;
	assert RAM(15110) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(15110))))  severity failure;
	assert RAM(15111) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15111))))  severity failure;
	assert RAM(15112) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(15112))))  severity failure;
	assert RAM(15113) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(15113))))  severity failure;
	assert RAM(15114) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(15114))))  severity failure;
	assert RAM(15115) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(15115))))  severity failure;
	assert RAM(15116) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(15116))))  severity failure;
	assert RAM(15117) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(15117))))  severity failure;
	assert RAM(15118) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(15118))))  severity failure;
	assert RAM(15119) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(15119))))  severity failure;
	assert RAM(15120) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(15120))))  severity failure;
	assert RAM(15121) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(15121))))  severity failure;
	assert RAM(15122) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(15122))))  severity failure;
	assert RAM(15123) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(15123))))  severity failure;
	assert RAM(15124) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(15124))))  severity failure;
	assert RAM(15125) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(15125))))  severity failure;
	assert RAM(15126) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(15126))))  severity failure;
	assert RAM(15127) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(15127))))  severity failure;
	assert RAM(15128) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(15128))))  severity failure;
	assert RAM(15129) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(15129))))  severity failure;
	assert RAM(15130) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(15130))))  severity failure;
	assert RAM(15131) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(15131))))  severity failure;
	assert RAM(15132) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(15132))))  severity failure;
	assert RAM(15133) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(15133))))  severity failure;
	assert RAM(15134) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(15134))))  severity failure;
	assert RAM(15135) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(15135))))  severity failure;
	assert RAM(15136) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(15136))))  severity failure;
	assert RAM(15137) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(15137))))  severity failure;
	assert RAM(15138) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(15138))))  severity failure;
	assert RAM(15139) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(15139))))  severity failure;
	assert RAM(15140) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(15140))))  severity failure;
	assert RAM(15141) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(15141))))  severity failure;
	assert RAM(15142) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15142))))  severity failure;
	assert RAM(15143) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(15143))))  severity failure;
	assert RAM(15144) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(15144))))  severity failure;
	assert RAM(15145) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(15145))))  severity failure;
	assert RAM(15146) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(15146))))  severity failure;
	assert RAM(15147) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(15147))))  severity failure;
	assert RAM(15148) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(15148))))  severity failure;
	assert RAM(15149) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(15149))))  severity failure;
	assert RAM(15150) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(15150))))  severity failure;
	assert RAM(15151) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(15151))))  severity failure;
	assert RAM(15152) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(15152))))  severity failure;
	assert RAM(15153) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(15153))))  severity failure;
	assert RAM(15154) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(15154))))  severity failure;
	assert RAM(15155) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(15155))))  severity failure;
	assert RAM(15156) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(15156))))  severity failure;
	assert RAM(15157) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(15157))))  severity failure;
	assert RAM(15158) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(15158))))  severity failure;
	assert RAM(15159) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(15159))))  severity failure;
	assert RAM(15160) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(15160))))  severity failure;
	assert RAM(15161) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(15161))))  severity failure;
	assert RAM(15162) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(15162))))  severity failure;
	assert RAM(15163) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(15163))))  severity failure;
	assert RAM(15164) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(15164))))  severity failure;
	assert RAM(15165) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(15165))))  severity failure;
	assert RAM(15166) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(15166))))  severity failure;
	assert RAM(15167) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(15167))))  severity failure;
	assert RAM(15168) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(15168))))  severity failure;
	assert RAM(15169) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15169))))  severity failure;
	assert RAM(15170) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(15170))))  severity failure;
	assert RAM(15171) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(15171))))  severity failure;
	assert RAM(15172) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(15172))))  severity failure;
	assert RAM(15173) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(15173))))  severity failure;
	assert RAM(15174) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(15174))))  severity failure;
	assert RAM(15175) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(15175))))  severity failure;
	assert RAM(15176) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(15176))))  severity failure;
	assert RAM(15177) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(15177))))  severity failure;
	assert RAM(15178) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(15178))))  severity failure;
	assert RAM(15179) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(15179))))  severity failure;
	assert RAM(15180) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(15180))))  severity failure;
	assert RAM(15181) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15181))))  severity failure;
	assert RAM(15182) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(15182))))  severity failure;
	assert RAM(15183) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(15183))))  severity failure;
	assert RAM(15184) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(15184))))  severity failure;
	assert RAM(15185) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(15185))))  severity failure;
	assert RAM(15186) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(15186))))  severity failure;
	assert RAM(15187) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(15187))))  severity failure;
	assert RAM(15188) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(15188))))  severity failure;
	assert RAM(15189) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(15189))))  severity failure;
	assert RAM(15190) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(15190))))  severity failure;
	assert RAM(15191) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(15191))))  severity failure;
	assert RAM(15192) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(15192))))  severity failure;
	assert RAM(15193) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(15193))))  severity failure;
	assert RAM(15194) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(15194))))  severity failure;
	assert RAM(15195) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(15195))))  severity failure;
	assert RAM(15196) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(15196))))  severity failure;
	assert RAM(15197) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(15197))))  severity failure;
	assert RAM(15198) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(15198))))  severity failure;
	assert RAM(15199) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(15199))))  severity failure;
	assert RAM(15200) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(15200))))  severity failure;
	assert RAM(15201) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(15201))))  severity failure;
	assert RAM(15202) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(15202))))  severity failure;
	assert RAM(15203) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(15203))))  severity failure;
	assert RAM(15204) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(15204))))  severity failure;
	assert RAM(15205) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(15205))))  severity failure;
	assert RAM(15206) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(15206))))  severity failure;
	assert RAM(15207) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(15207))))  severity failure;
	assert RAM(15208) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(15208))))  severity failure;
	assert RAM(15209) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(15209))))  severity failure;
	assert RAM(15210) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(15210))))  severity failure;
	assert RAM(15211) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(15211))))  severity failure;
	assert RAM(15212) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(15212))))  severity failure;
	assert RAM(15213) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(15213))))  severity failure;
	assert RAM(15214) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(15214))))  severity failure;
	assert RAM(15215) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(15215))))  severity failure;
	assert RAM(15216) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(15216))))  severity failure;
	assert RAM(15217) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(15217))))  severity failure;
	assert RAM(15218) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(15218))))  severity failure;
	assert RAM(15219) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(15219))))  severity failure;
	assert RAM(15220) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15220))))  severity failure;
	assert RAM(15221) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(15221))))  severity failure;
	assert RAM(15222) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(15222))))  severity failure;
	assert RAM(15223) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(15223))))  severity failure;
	assert RAM(15224) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(15224))))  severity failure;
	assert RAM(15225) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(15225))))  severity failure;
	assert RAM(15226) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(15226))))  severity failure;
	assert RAM(15227) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15227))))  severity failure;
	assert RAM(15228) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(15228))))  severity failure;
	assert RAM(15229) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(15229))))  severity failure;
	assert RAM(15230) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(15230))))  severity failure;
	assert RAM(15231) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(15231))))  severity failure;
	assert RAM(15232) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(15232))))  severity failure;
	assert RAM(15233) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15233))))  severity failure;
	assert RAM(15234) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(15234))))  severity failure;
	assert RAM(15235) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(15235))))  severity failure;
	assert RAM(15236) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(15236))))  severity failure;
	assert RAM(15237) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(15237))))  severity failure;
	assert RAM(15238) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(15238))))  severity failure;
	assert RAM(15239) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(15239))))  severity failure;
	assert RAM(15240) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(15240))))  severity failure;
	assert RAM(15241) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(15241))))  severity failure;
	assert RAM(15242) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15242))))  severity failure;
	assert RAM(15243) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(15243))))  severity failure;
	assert RAM(15244) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(15244))))  severity failure;
	assert RAM(15245) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(15245))))  severity failure;
	assert RAM(15246) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(15246))))  severity failure;
	assert RAM(15247) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(15247))))  severity failure;
	assert RAM(15248) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(15248))))  severity failure;
	assert RAM(15249) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(15249))))  severity failure;
	assert RAM(15250) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(15250))))  severity failure;
	assert RAM(15251) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(15251))))  severity failure;
	assert RAM(15252) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(15252))))  severity failure;
	assert RAM(15253) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(15253))))  severity failure;
	assert RAM(15254) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(15254))))  severity failure;
	assert RAM(15255) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(15255))))  severity failure;
	assert RAM(15256) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(15256))))  severity failure;
	assert RAM(15257) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(15257))))  severity failure;
	assert RAM(15258) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(15258))))  severity failure;
	assert RAM(15259) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(15259))))  severity failure;
	assert RAM(15260) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(15260))))  severity failure;
	assert RAM(15261) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(15261))))  severity failure;
	assert RAM(15262) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(15262))))  severity failure;
	assert RAM(15263) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(15263))))  severity failure;
	assert RAM(15264) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(15264))))  severity failure;
	assert RAM(15265) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(15265))))  severity failure;
	assert RAM(15266) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(15266))))  severity failure;
	assert RAM(15267) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(15267))))  severity failure;
	assert RAM(15268) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(15268))))  severity failure;
	assert RAM(15269) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(15269))))  severity failure;
	assert RAM(15270) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(15270))))  severity failure;
	assert RAM(15271) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(15271))))  severity failure;
	assert RAM(15272) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(15272))))  severity failure;
	assert RAM(15273) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(15273))))  severity failure;
	assert RAM(15274) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(15274))))  severity failure;
	assert RAM(15275) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(15275))))  severity failure;
	assert RAM(15276) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(15276))))  severity failure;
	assert RAM(15277) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(15277))))  severity failure;
	assert RAM(15278) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(15278))))  severity failure;
	assert RAM(15279) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(15279))))  severity failure;
	assert RAM(15280) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(15280))))  severity failure;
	assert RAM(15281) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(15281))))  severity failure;
	assert RAM(15282) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(15282))))  severity failure;
	assert RAM(15283) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(15283))))  severity failure;
	assert RAM(15284) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(15284))))  severity failure;
	assert RAM(15285) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(15285))))  severity failure;
	assert RAM(15286) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(15286))))  severity failure;
	assert RAM(15287) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(15287))))  severity failure;
	assert RAM(15288) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(15288))))  severity failure;
	assert RAM(15289) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(15289))))  severity failure;
	assert RAM(15290) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(15290))))  severity failure;
	assert RAM(15291) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(15291))))  severity failure;
	assert RAM(15292) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(15292))))  severity failure;
	assert RAM(15293) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(15293))))  severity failure;
	assert RAM(15294) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(15294))))  severity failure;
	assert RAM(15295) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(15295))))  severity failure;
	assert RAM(15296) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(15296))))  severity failure;
	assert RAM(15297) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(15297))))  severity failure;
	assert RAM(15298) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(15298))))  severity failure;
	assert RAM(15299) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(15299))))  severity failure;
	assert RAM(15300) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(15300))))  severity failure;
	assert RAM(15301) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(15301))))  severity failure;
	assert RAM(15302) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(15302))))  severity failure;
	assert RAM(15303) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(15303))))  severity failure;
	assert RAM(15304) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(15304))))  severity failure;
	assert RAM(15305) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(15305))))  severity failure;
	assert RAM(15306) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(15306))))  severity failure;
	assert RAM(15307) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(15307))))  severity failure;
	assert RAM(15308) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(15308))))  severity failure;
	assert RAM(15309) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(15309))))  severity failure;
	assert RAM(15310) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(15310))))  severity failure;
	assert RAM(15311) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(15311))))  severity failure;
	assert RAM(15312) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(15312))))  severity failure;
	assert RAM(15313) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(15313))))  severity failure;
	assert RAM(15314) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(15314))))  severity failure;
	assert RAM(15315) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(15315))))  severity failure;
	assert RAM(15316) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(15316))))  severity failure;
	assert RAM(15317) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15317))))  severity failure;
	assert RAM(15318) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(15318))))  severity failure;
	assert RAM(15319) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(15319))))  severity failure;
	assert RAM(15320) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(15320))))  severity failure;
	assert RAM(15321) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(15321))))  severity failure;
	assert RAM(15322) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(15322))))  severity failure;
	assert RAM(15323) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(15323))))  severity failure;
	assert RAM(15324) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(15324))))  severity failure;
	assert RAM(15325) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(15325))))  severity failure;
	assert RAM(15326) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(15326))))  severity failure;
	assert RAM(15327) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(15327))))  severity failure;
	assert RAM(15328) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(15328))))  severity failure;
	assert RAM(15329) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(15329))))  severity failure;
	assert RAM(15330) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(15330))))  severity failure;
	assert RAM(15331) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(15331))))  severity failure;
	assert RAM(15332) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15332))))  severity failure;
	assert RAM(15333) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(15333))))  severity failure;
	assert RAM(15334) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(15334))))  severity failure;
	assert RAM(15335) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(15335))))  severity failure;
	assert RAM(15336) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(15336))))  severity failure;
	assert RAM(15337) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(15337))))  severity failure;
	assert RAM(15338) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(15338))))  severity failure;
	assert RAM(15339) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(15339))))  severity failure;
	assert RAM(15340) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(15340))))  severity failure;
	assert RAM(15341) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(15341))))  severity failure;
	assert RAM(15342) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(15342))))  severity failure;
	assert RAM(15343) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(15343))))  severity failure;
	assert RAM(15344) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(15344))))  severity failure;
	assert RAM(15345) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(15345))))  severity failure;
	assert RAM(15346) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(15346))))  severity failure;
	assert RAM(15347) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(15347))))  severity failure;
	assert RAM(15348) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(15348))))  severity failure;
	assert RAM(15349) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(15349))))  severity failure;
	assert RAM(15350) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(15350))))  severity failure;
	assert RAM(15351) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(15351))))  severity failure;
	assert RAM(15352) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(15352))))  severity failure;
	assert RAM(15353) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(15353))))  severity failure;
	assert RAM(15354) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(15354))))  severity failure;
	assert RAM(15355) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(15355))))  severity failure;
	assert RAM(15356) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(15356))))  severity failure;
	assert RAM(15357) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(15357))))  severity failure;
	assert RAM(15358) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(15358))))  severity failure;
	assert RAM(15359) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(15359))))  severity failure;
	assert RAM(15360) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(15360))))  severity failure;
	assert RAM(15361) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(15361))))  severity failure;
	assert RAM(15362) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(15362))))  severity failure;
	assert RAM(15363) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(15363))))  severity failure;
	assert RAM(15364) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(15364))))  severity failure;
	assert RAM(15365) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(15365))))  severity failure;
	assert RAM(15366) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(15366))))  severity failure;
	assert RAM(15367) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(15367))))  severity failure;
	assert RAM(15368) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(15368))))  severity failure;
	assert RAM(15369) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(15369))))  severity failure;
	assert RAM(15370) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(15370))))  severity failure;
	assert RAM(15371) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(15371))))  severity failure;
	assert RAM(15372) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(15372))))  severity failure;
	assert RAM(15373) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(15373))))  severity failure;
	assert RAM(15374) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(15374))))  severity failure;
	assert RAM(15375) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(15375))))  severity failure;
	assert RAM(15376) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(15376))))  severity failure;
	assert RAM(15377) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(15377))))  severity failure;
	assert RAM(15378) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(15378))))  severity failure;
	assert RAM(15379) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(15379))))  severity failure;
	assert RAM(15380) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(15380))))  severity failure;
	assert RAM(15381) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(15381))))  severity failure;
	assert RAM(15382) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(15382))))  severity failure;
	assert RAM(15383) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(15383))))  severity failure;
	assert RAM(15384) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(15384))))  severity failure;
	assert RAM(15385) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(15385))))  severity failure;
	assert RAM(15386) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(15386))))  severity failure;
	assert RAM(15387) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(15387))))  severity failure;
	assert RAM(15388) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(15388))))  severity failure;
	assert RAM(15389) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(15389))))  severity failure;
	assert RAM(15390) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(15390))))  severity failure;
	assert RAM(15391) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(15391))))  severity failure;
	assert RAM(15392) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(15392))))  severity failure;
	assert RAM(15393) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(15393))))  severity failure;
	assert RAM(15394) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(15394))))  severity failure;
	assert RAM(15395) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(15395))))  severity failure;
	assert RAM(15396) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(15396))))  severity failure;
	assert RAM(15397) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(15397))))  severity failure;
	assert RAM(15398) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(15398))))  severity failure;
	assert RAM(15399) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(15399))))  severity failure;
	assert RAM(15400) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(15400))))  severity failure;
	assert RAM(15401) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(15401))))  severity failure;
	assert RAM(15402) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(15402))))  severity failure;
	assert RAM(15403) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(15403))))  severity failure;
	assert RAM(15404) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(15404))))  severity failure;
	assert RAM(15405) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(15405))))  severity failure;
	assert RAM(15406) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15406))))  severity failure;
	assert RAM(15407) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(15407))))  severity failure;
	assert RAM(15408) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(15408))))  severity failure;
	assert RAM(15409) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15409))))  severity failure;
	assert RAM(15410) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(15410))))  severity failure;
	assert RAM(15411) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(15411))))  severity failure;
	assert RAM(15412) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(15412))))  severity failure;
	assert RAM(15413) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(15413))))  severity failure;
	assert RAM(15414) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(15414))))  severity failure;
	assert RAM(15415) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(15415))))  severity failure;
	assert RAM(15416) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(15416))))  severity failure;
	assert RAM(15417) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(15417))))  severity failure;
	assert RAM(15418) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(15418))))  severity failure;
	assert RAM(15419) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(15419))))  severity failure;
	assert RAM(15420) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(15420))))  severity failure;
	assert RAM(15421) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(15421))))  severity failure;
	assert RAM(15422) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(15422))))  severity failure;
	assert RAM(15423) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(15423))))  severity failure;
	assert RAM(15424) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(15424))))  severity failure;
	assert RAM(15425) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(15425))))  severity failure;
	assert RAM(15426) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(15426))))  severity failure;
	assert RAM(15427) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(15427))))  severity failure;
	assert RAM(15428) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(15428))))  severity failure;
	assert RAM(15429) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(15429))))  severity failure;
	assert RAM(15430) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(15430))))  severity failure;
	assert RAM(15431) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(15431))))  severity failure;
	assert RAM(15432) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(15432))))  severity failure;
	assert RAM(15433) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(15433))))  severity failure;
	assert RAM(15434) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(15434))))  severity failure;
	assert RAM(15435) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(15435))))  severity failure;
	assert RAM(15436) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(15436))))  severity failure;
	assert RAM(15437) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(15437))))  severity failure;
	assert RAM(15438) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(15438))))  severity failure;
	assert RAM(15439) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(15439))))  severity failure;
	assert RAM(15440) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(15440))))  severity failure;
	assert RAM(15441) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(15441))))  severity failure;
	assert RAM(15442) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(15442))))  severity failure;
	assert RAM(15443) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(15443))))  severity failure;
	assert RAM(15444) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(15444))))  severity failure;
	assert RAM(15445) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(15445))))  severity failure;
	assert RAM(15446) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(15446))))  severity failure;
	assert RAM(15447) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(15447))))  severity failure;
	assert RAM(15448) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(15448))))  severity failure;
	assert RAM(15449) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(15449))))  severity failure;
	assert RAM(15450) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(15450))))  severity failure;
	assert RAM(15451) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(15451))))  severity failure;
	assert RAM(15452) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(15452))))  severity failure;
	assert RAM(15453) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(15453))))  severity failure;
	assert RAM(15454) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(15454))))  severity failure;
	assert RAM(15455) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(15455))))  severity failure;
	assert RAM(15456) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(15456))))  severity failure;
	assert RAM(15457) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(15457))))  severity failure;
	assert RAM(15458) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(15458))))  severity failure;
	assert RAM(15459) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(15459))))  severity failure;
	assert RAM(15460) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(15460))))  severity failure;
	assert RAM(15461) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(15461))))  severity failure;
	assert RAM(15462) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(15462))))  severity failure;
	assert RAM(15463) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(15463))))  severity failure;
	assert RAM(15464) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(15464))))  severity failure;
	assert RAM(15465) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(15465))))  severity failure;
	assert RAM(15466) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(15466))))  severity failure;
	assert RAM(15467) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(15467))))  severity failure;
	assert RAM(15468) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(15468))))  severity failure;
	assert RAM(15469) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(15469))))  severity failure;
	assert RAM(15470) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(15470))))  severity failure;
	assert RAM(15471) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(15471))))  severity failure;
	assert RAM(15472) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(15472))))  severity failure;
	assert RAM(15473) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(15473))))  severity failure;
	assert RAM(15474) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(15474))))  severity failure;
	assert RAM(15475) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(15475))))  severity failure;
	assert RAM(15476) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(15476))))  severity failure;
	assert RAM(15477) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(15477))))  severity failure;
	assert RAM(15478) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(15478))))  severity failure;
	assert RAM(15479) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(15479))))  severity failure;
	assert RAM(15480) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(15480))))  severity failure;
	assert RAM(15481) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(15481))))  severity failure;
	assert RAM(15482) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(15482))))  severity failure;
	assert RAM(15483) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(15483))))  severity failure;
	assert RAM(15484) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(15484))))  severity failure;
	assert RAM(15485) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(15485))))  severity failure;
	assert RAM(15486) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(15486))))  severity failure;
	assert RAM(15487) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(15487))))  severity failure;
	assert RAM(15488) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15488))))  severity failure;
	assert RAM(15489) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(15489))))  severity failure;
	assert RAM(15490) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(15490))))  severity failure;
	assert RAM(15491) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(15491))))  severity failure;
	assert RAM(15492) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(15492))))  severity failure;
	assert RAM(15493) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(15493))))  severity failure;
	assert RAM(15494) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(15494))))  severity failure;
	assert RAM(15495) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(15495))))  severity failure;
	assert RAM(15496) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(15496))))  severity failure;
	assert RAM(15497) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(15497))))  severity failure;
	assert RAM(15498) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(15498))))  severity failure;
	assert RAM(15499) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(15499))))  severity failure;
	assert RAM(15500) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(15500))))  severity failure;
	assert RAM(15501) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(15501))))  severity failure;
	assert RAM(15502) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(15502))))  severity failure;
	assert RAM(15503) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(15503))))  severity failure;
	assert RAM(15504) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(15504))))  severity failure;
	assert RAM(15505) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(15505))))  severity failure;
	assert RAM(15506) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(15506))))  severity failure;
	assert RAM(15507) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(15507))))  severity failure;
	assert RAM(15508) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(15508))))  severity failure;
	assert RAM(15509) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(15509))))  severity failure;
	assert RAM(15510) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(15510))))  severity failure;
	assert RAM(15511) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(15511))))  severity failure;
	assert RAM(15512) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15512))))  severity failure;
	assert RAM(15513) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(15513))))  severity failure;
	assert RAM(15514) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(15514))))  severity failure;
	assert RAM(15515) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(15515))))  severity failure;
	assert RAM(15516) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(15516))))  severity failure;
	assert RAM(15517) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(15517))))  severity failure;
	assert RAM(15518) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(15518))))  severity failure;
	assert RAM(15519) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(15519))))  severity failure;
	assert RAM(15520) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(15520))))  severity failure;
	assert RAM(15521) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(15521))))  severity failure;
	assert RAM(15522) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(15522))))  severity failure;
	assert RAM(15523) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(15523))))  severity failure;
	assert RAM(15524) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(15524))))  severity failure;
	assert RAM(15525) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(15525))))  severity failure;
	assert RAM(15526) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(15526))))  severity failure;
	assert RAM(15527) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(15527))))  severity failure;
	assert RAM(15528) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(15528))))  severity failure;
	assert RAM(15529) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(15529))))  severity failure;
	assert RAM(15530) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(15530))))  severity failure;
	assert RAM(15531) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(15531))))  severity failure;
	assert RAM(15532) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(15532))))  severity failure;
	assert RAM(15533) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(15533))))  severity failure;
	assert RAM(15534) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(15534))))  severity failure;
	assert RAM(15535) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(15535))))  severity failure;
	assert RAM(15536) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(15536))))  severity failure;
	assert RAM(15537) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(15537))))  severity failure;
	assert RAM(15538) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(15538))))  severity failure;
	assert RAM(15539) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(15539))))  severity failure;
	assert RAM(15540) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(15540))))  severity failure;
	assert RAM(15541) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(15541))))  severity failure;
	assert RAM(15542) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(15542))))  severity failure;
	assert RAM(15543) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(15543))))  severity failure;
	assert RAM(15544) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(15544))))  severity failure;
	assert RAM(15545) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(15545))))  severity failure;
	assert RAM(15546) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(15546))))  severity failure;
	assert RAM(15547) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(15547))))  severity failure;
	assert RAM(15548) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(15548))))  severity failure;
	assert RAM(15549) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(15549))))  severity failure;
	assert RAM(15550) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(15550))))  severity failure;
	assert RAM(15551) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(15551))))  severity failure;
	assert RAM(15552) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(15552))))  severity failure;
	assert RAM(15553) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(15553))))  severity failure;
	assert RAM(15554) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15554))))  severity failure;
	assert RAM(15555) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(15555))))  severity failure;
	assert RAM(15556) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(15556))))  severity failure;
	assert RAM(15557) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15557))))  severity failure;
	assert RAM(15558) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(15558))))  severity failure;
	assert RAM(15559) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(15559))))  severity failure;
	assert RAM(15560) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(15560))))  severity failure;
	assert RAM(15561) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(15561))))  severity failure;
	assert RAM(15562) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(15562))))  severity failure;
	assert RAM(15563) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(15563))))  severity failure;
	assert RAM(15564) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(15564))))  severity failure;
	assert RAM(15565) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(15565))))  severity failure;
	assert RAM(15566) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(15566))))  severity failure;
	assert RAM(15567) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(15567))))  severity failure;
	assert RAM(15568) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(15568))))  severity failure;
	assert RAM(15569) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(15569))))  severity failure;
	assert RAM(15570) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(15570))))  severity failure;
	assert RAM(15571) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15571))))  severity failure;
	assert RAM(15572) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(15572))))  severity failure;
	assert RAM(15573) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(15573))))  severity failure;
	assert RAM(15574) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(15574))))  severity failure;
	assert RAM(15575) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(15575))))  severity failure;
	assert RAM(15576) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(15576))))  severity failure;
	assert RAM(15577) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(15577))))  severity failure;
	assert RAM(15578) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(15578))))  severity failure;
	assert RAM(15579) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(15579))))  severity failure;
	assert RAM(15580) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(15580))))  severity failure;
	assert RAM(15581) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15581))))  severity failure;
	assert RAM(15582) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(15582))))  severity failure;
	assert RAM(15583) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(15583))))  severity failure;
	assert RAM(15584) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(15584))))  severity failure;
	assert RAM(15585) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(15585))))  severity failure;
	assert RAM(15586) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(15586))))  severity failure;
	assert RAM(15587) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(15587))))  severity failure;
	assert RAM(15588) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(15588))))  severity failure;
	assert RAM(15589) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(15589))))  severity failure;
	assert RAM(15590) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(15590))))  severity failure;
	assert RAM(15591) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(15591))))  severity failure;
	assert RAM(15592) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(15592))))  severity failure;
	assert RAM(15593) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(15593))))  severity failure;
	assert RAM(15594) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(15594))))  severity failure;
	assert RAM(15595) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(15595))))  severity failure;
	assert RAM(15596) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(15596))))  severity failure;
	assert RAM(15597) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(15597))))  severity failure;
	assert RAM(15598) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(15598))))  severity failure;
	assert RAM(15599) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(15599))))  severity failure;
	assert RAM(15600) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(15600))))  severity failure;
	assert RAM(15601) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(15601))))  severity failure;
	assert RAM(15602) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(15602))))  severity failure;
	assert RAM(15603) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(15603))))  severity failure;
	assert RAM(15604) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(15604))))  severity failure;
	assert RAM(15605) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(15605))))  severity failure;
	assert RAM(15606) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(15606))))  severity failure;
	assert RAM(15607) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(15607))))  severity failure;
	assert RAM(15608) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(15608))))  severity failure;
	assert RAM(15609) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(15609))))  severity failure;
	assert RAM(15610) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(15610))))  severity failure;
	assert RAM(15611) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(15611))))  severity failure;
	assert RAM(15612) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(15612))))  severity failure;
	assert RAM(15613) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(15613))))  severity failure;
	assert RAM(15614) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(15614))))  severity failure;
	assert RAM(15615) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(15615))))  severity failure;
	assert RAM(15616) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(15616))))  severity failure;
	assert RAM(15617) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(15617))))  severity failure;
	assert RAM(15618) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(15618))))  severity failure;
	assert RAM(15619) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(15619))))  severity failure;
	assert RAM(15620) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(15620))))  severity failure;
	assert RAM(15621) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(15621))))  severity failure;
	assert RAM(15622) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(15622))))  severity failure;
	assert RAM(15623) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(15623))))  severity failure;
	assert RAM(15624) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(15624))))  severity failure;
	assert RAM(15625) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(15625))))  severity failure;
	assert RAM(15626) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(15626))))  severity failure;
	assert RAM(15627) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(15627))))  severity failure;
	assert RAM(15628) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(15628))))  severity failure;
	assert RAM(15629) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(15629))))  severity failure;
	assert RAM(15630) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(15630))))  severity failure;
	assert RAM(15631) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(15631))))  severity failure;
	assert RAM(15632) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(15632))))  severity failure;
	assert RAM(15633) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(15633))))  severity failure;
	assert RAM(15634) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(15634))))  severity failure;
	assert RAM(15635) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(15635))))  severity failure;
	assert RAM(15636) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(15636))))  severity failure;
	assert RAM(15637) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(15637))))  severity failure;
	assert RAM(15638) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(15638))))  severity failure;
	assert RAM(15639) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(15639))))  severity failure;
	assert RAM(15640) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(15640))))  severity failure;
	assert RAM(15641) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(15641))))  severity failure;
	assert RAM(15642) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(15642))))  severity failure;
	assert RAM(15643) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(15643))))  severity failure;
	assert RAM(15644) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(15644))))  severity failure;
	assert RAM(15645) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(15645))))  severity failure;
	assert RAM(15646) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(15646))))  severity failure;
	assert RAM(15647) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(15647))))  severity failure;
	assert RAM(15648) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(15648))))  severity failure;
	assert RAM(15649) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(15649))))  severity failure;
	assert RAM(15650) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(15650))))  severity failure;
	assert RAM(15651) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(15651))))  severity failure;
	assert RAM(15652) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(15652))))  severity failure;
	assert RAM(15653) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(15653))))  severity failure;
	assert RAM(15654) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(15654))))  severity failure;
	assert RAM(15655) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(15655))))  severity failure;
	assert RAM(15656) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(15656))))  severity failure;
	assert RAM(15657) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(15657))))  severity failure;
	assert RAM(15658) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(15658))))  severity failure;
	assert RAM(15659) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(15659))))  severity failure;
	assert RAM(15660) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(15660))))  severity failure;
	assert RAM(15661) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(15661))))  severity failure;
	assert RAM(15662) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(15662))))  severity failure;
	assert RAM(15663) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(15663))))  severity failure;
	assert RAM(15664) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(15664))))  severity failure;
	assert RAM(15665) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(15665))))  severity failure;
	assert RAM(15666) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(15666))))  severity failure;
	assert RAM(15667) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(15667))))  severity failure;
	assert RAM(15668) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(15668))))  severity failure;
	assert RAM(15669) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(15669))))  severity failure;
	assert RAM(15670) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(15670))))  severity failure;
	assert RAM(15671) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(15671))))  severity failure;
	assert RAM(15672) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(15672))))  severity failure;
	assert RAM(15673) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(15673))))  severity failure;
	assert RAM(15674) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(15674))))  severity failure;
	assert RAM(15675) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(15675))))  severity failure;
	assert RAM(15676) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(15676))))  severity failure;
	assert RAM(15677) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(15677))))  severity failure;
	assert RAM(15678) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(15678))))  severity failure;
	assert RAM(15679) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(15679))))  severity failure;
	assert RAM(15680) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(15680))))  severity failure;
	assert RAM(15681) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(15681))))  severity failure;
	assert RAM(15682) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(15682))))  severity failure;
	assert RAM(15683) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(15683))))  severity failure;
	assert RAM(15684) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(15684))))  severity failure;
	assert RAM(15685) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(15685))))  severity failure;
	assert RAM(15686) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(15686))))  severity failure;
	assert RAM(15687) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(15687))))  severity failure;
	assert RAM(15688) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(15688))))  severity failure;
	assert RAM(15689) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(15689))))  severity failure;
	assert RAM(15690) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(15690))))  severity failure;
	assert RAM(15691) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(15691))))  severity failure;
	assert RAM(15692) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(15692))))  severity failure;
	assert RAM(15693) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(15693))))  severity failure;
	assert RAM(15694) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(15694))))  severity failure;
	assert RAM(15695) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(15695))))  severity failure;
	assert RAM(15696) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(15696))))  severity failure;
	assert RAM(15697) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(15697))))  severity failure;
	assert RAM(15698) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(15698))))  severity failure;
	assert RAM(15699) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(15699))))  severity failure;
	assert RAM(15700) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(15700))))  severity failure;
	assert RAM(15701) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(15701))))  severity failure;
	assert RAM(15702) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(15702))))  severity failure;
	assert RAM(15703) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(15703))))  severity failure;
	assert RAM(15704) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(15704))))  severity failure;
	assert RAM(15705) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(15705))))  severity failure;
	assert RAM(15706) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(15706))))  severity failure;
	assert RAM(15707) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(15707))))  severity failure;
	assert RAM(15708) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(15708))))  severity failure;
	assert RAM(15709) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(15709))))  severity failure;
	assert RAM(15710) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(15710))))  severity failure;
	assert RAM(15711) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(15711))))  severity failure;
	assert RAM(15712) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(15712))))  severity failure;
	assert RAM(15713) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(15713))))  severity failure;
	assert RAM(15714) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(15714))))  severity failure;
	assert RAM(15715) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(15715))))  severity failure;
	assert RAM(15716) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(15716))))  severity failure;
	assert RAM(15717) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(15717))))  severity failure;
	assert RAM(15718) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(15718))))  severity failure;
	assert RAM(15719) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(15719))))  severity failure;
	assert RAM(15720) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(15720))))  severity failure;
	assert RAM(15721) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(15721))))  severity failure;
	assert RAM(15722) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(15722))))  severity failure;
	assert RAM(15723) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(15723))))  severity failure;
	assert RAM(15724) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(15724))))  severity failure;
	assert RAM(15725) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(15725))))  severity failure;
	assert RAM(15726) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(15726))))  severity failure;
	assert RAM(15727) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(15727))))  severity failure;
	assert RAM(15728) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(15728))))  severity failure;
	assert RAM(15729) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(15729))))  severity failure;
	assert RAM(15730) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(15730))))  severity failure;
	assert RAM(15731) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(15731))))  severity failure;
	assert RAM(15732) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(15732))))  severity failure;
	assert RAM(15733) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(15733))))  severity failure;
	assert RAM(15734) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(15734))))  severity failure;
	assert RAM(15735) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(15735))))  severity failure;
	assert RAM(15736) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(15736))))  severity failure;
	assert RAM(15737) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(15737))))  severity failure;
	assert RAM(15738) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(15738))))  severity failure;
	assert RAM(15739) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(15739))))  severity failure;
	assert RAM(15740) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(15740))))  severity failure;
	assert RAM(15741) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(15741))))  severity failure;
	assert RAM(15742) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(15742))))  severity failure;
	assert RAM(15743) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(15743))))  severity failure;
	assert RAM(15744) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(15744))))  severity failure;
	assert RAM(15745) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(15745))))  severity failure;
	assert RAM(15746) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15746))))  severity failure;
	assert RAM(15747) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(15747))))  severity failure;
	assert RAM(15748) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(15748))))  severity failure;
	assert RAM(15749) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(15749))))  severity failure;
	assert RAM(15750) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(15750))))  severity failure;
	assert RAM(15751) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(15751))))  severity failure;
	assert RAM(15752) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(15752))))  severity failure;
	assert RAM(15753) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(15753))))  severity failure;
	assert RAM(15754) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(15754))))  severity failure;
	assert RAM(15755) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(15755))))  severity failure;
	assert RAM(15756) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(15756))))  severity failure;
	assert RAM(15757) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(15757))))  severity failure;
	assert RAM(15758) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(15758))))  severity failure;
	assert RAM(15759) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(15759))))  severity failure;
	assert RAM(15760) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(15760))))  severity failure;
	assert RAM(15761) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(15761))))  severity failure;
	assert RAM(15762) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(15762))))  severity failure;
	assert RAM(15763) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(15763))))  severity failure;
	assert RAM(15764) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(15764))))  severity failure;
	assert RAM(15765) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(15765))))  severity failure;
	assert RAM(15766) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(15766))))  severity failure;
	assert RAM(15767) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(15767))))  severity failure;
	assert RAM(15768) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(15768))))  severity failure;
	assert RAM(15769) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(15769))))  severity failure;
	assert RAM(15770) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(15770))))  severity failure;
	assert RAM(15771) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(15771))))  severity failure;
	assert RAM(15772) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(15772))))  severity failure;
	assert RAM(15773) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(15773))))  severity failure;
	assert RAM(15774) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(15774))))  severity failure;
	assert RAM(15775) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(15775))))  severity failure;
	assert RAM(15776) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(15776))))  severity failure;
	assert RAM(15777) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(15777))))  severity failure;
	assert RAM(15778) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(15778))))  severity failure;
	assert RAM(15779) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(15779))))  severity failure;
	assert RAM(15780) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(15780))))  severity failure;
	assert RAM(15781) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(15781))))  severity failure;
	assert RAM(15782) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(15782))))  severity failure;
	assert RAM(15783) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(15783))))  severity failure;
	assert RAM(15784) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(15784))))  severity failure;
	assert RAM(15785) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(15785))))  severity failure;
	assert RAM(15786) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(15786))))  severity failure;
	assert RAM(15787) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(15787))))  severity failure;
	assert RAM(15788) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(15788))))  severity failure;
	assert RAM(15789) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(15789))))  severity failure;
	assert RAM(15790) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(15790))))  severity failure;
	assert RAM(15791) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(15791))))  severity failure;
	assert RAM(15792) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(15792))))  severity failure;
	assert RAM(15793) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(15793))))  severity failure;
	assert RAM(15794) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(15794))))  severity failure;
	assert RAM(15795) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(15795))))  severity failure;
	assert RAM(15796) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(15796))))  severity failure;
	assert RAM(15797) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(15797))))  severity failure;
	assert RAM(15798) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(15798))))  severity failure;
	assert RAM(15799) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(15799))))  severity failure;
	assert RAM(15800) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(15800))))  severity failure;
	assert RAM(15801) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(15801))))  severity failure;
	assert RAM(15802) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(15802))))  severity failure;
	assert RAM(15803) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(15803))))  severity failure;
	assert RAM(15804) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(15804))))  severity failure;
	assert RAM(15805) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(15805))))  severity failure;
	assert RAM(15806) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(15806))))  severity failure;
	assert RAM(15807) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(15807))))  severity failure;
	assert RAM(15808) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(15808))))  severity failure;
	assert RAM(15809) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(15809))))  severity failure;
	assert RAM(15810) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(15810))))  severity failure;
	assert RAM(15811) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(15811))))  severity failure;
	assert RAM(15812) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(15812))))  severity failure;
	assert RAM(15813) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(15813))))  severity failure;
	assert RAM(15814) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(15814))))  severity failure;
	assert RAM(15815) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(15815))))  severity failure;
	assert RAM(15816) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(15816))))  severity failure;
	assert RAM(15817) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(15817))))  severity failure;
	assert RAM(15818) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(15818))))  severity failure;
	assert RAM(15819) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(15819))))  severity failure;
	assert RAM(15820) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(15820))))  severity failure;
	assert RAM(15821) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(15821))))  severity failure;
	assert RAM(15822) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(15822))))  severity failure;
	assert RAM(15823) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(15823))))  severity failure;
	assert RAM(15824) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(15824))))  severity failure;
	assert RAM(15825) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(15825))))  severity failure;
	assert RAM(15826) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(15826))))  severity failure;
	assert RAM(15827) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(15827))))  severity failure;
	assert RAM(15828) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(15828))))  severity failure;
	assert RAM(15829) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(15829))))  severity failure;
	assert RAM(15830) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(15830))))  severity failure;
	assert RAM(15831) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(15831))))  severity failure;
	assert RAM(15832) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(15832))))  severity failure;
	assert RAM(15833) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(15833))))  severity failure;
	assert RAM(15834) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(15834))))  severity failure;
	assert RAM(15835) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(15835))))  severity failure;
	assert RAM(15836) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(15836))))  severity failure;
	assert RAM(15837) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(15837))))  severity failure;
	assert RAM(15838) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(15838))))  severity failure;
	assert RAM(15839) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(15839))))  severity failure;
	assert RAM(15840) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(15840))))  severity failure;
	assert RAM(15841) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(15841))))  severity failure;
	assert RAM(15842) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(15842))))  severity failure;
	assert RAM(15843) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(15843))))  severity failure;
	assert RAM(15844) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(15844))))  severity failure;
	assert RAM(15845) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(15845))))  severity failure;
	assert RAM(15846) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(15846))))  severity failure;
	assert RAM(15847) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(15847))))  severity failure;
	assert RAM(15848) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(15848))))  severity failure;
	assert RAM(15849) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(15849))))  severity failure;
	assert RAM(15850) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(15850))))  severity failure;
	assert RAM(15851) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15851))))  severity failure;
	assert RAM(15852) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(15852))))  severity failure;
	assert RAM(15853) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(15853))))  severity failure;
	assert RAM(15854) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(15854))))  severity failure;
	assert RAM(15855) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(15855))))  severity failure;
	assert RAM(15856) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(15856))))  severity failure;
	assert RAM(15857) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(15857))))  severity failure;
	assert RAM(15858) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(15858))))  severity failure;
	assert RAM(15859) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(15859))))  severity failure;
	assert RAM(15860) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(15860))))  severity failure;
	assert RAM(15861) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(15861))))  severity failure;
	assert RAM(15862) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(15862))))  severity failure;
	assert RAM(15863) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(15863))))  severity failure;
	assert RAM(15864) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(15864))))  severity failure;
	assert RAM(15865) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(15865))))  severity failure;
	assert RAM(15866) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(15866))))  severity failure;
	assert RAM(15867) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(15867))))  severity failure;
	assert RAM(15868) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(15868))))  severity failure;
	assert RAM(15869) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(15869))))  severity failure;
	assert RAM(15870) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(15870))))  severity failure;
	assert RAM(15871) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(15871))))  severity failure;
	assert RAM(15872) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(15872))))  severity failure;
	assert RAM(15873) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(15873))))  severity failure;
	assert RAM(15874) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(15874))))  severity failure;
	assert RAM(15875) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(15875))))  severity failure;
	assert RAM(15876) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(15876))))  severity failure;
	assert RAM(15877) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(15877))))  severity failure;
	assert RAM(15878) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(15878))))  severity failure;
	assert RAM(15879) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(15879))))  severity failure;
	assert RAM(15880) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(15880))))  severity failure;
	assert RAM(15881) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(15881))))  severity failure;
	assert RAM(15882) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(15882))))  severity failure;
	assert RAM(15883) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(15883))))  severity failure;
	assert RAM(15884) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(15884))))  severity failure;
	assert RAM(15885) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(15885))))  severity failure;
	assert RAM(15886) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(15886))))  severity failure;
	assert RAM(15887) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(15887))))  severity failure;
	assert RAM(15888) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(15888))))  severity failure;
	assert RAM(15889) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(15889))))  severity failure;
	assert RAM(15890) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(15890))))  severity failure;
	assert RAM(15891) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(15891))))  severity failure;
	assert RAM(15892) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(15892))))  severity failure;
	assert RAM(15893) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(15893))))  severity failure;
	assert RAM(15894) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(15894))))  severity failure;
	assert RAM(15895) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(15895))))  severity failure;
	assert RAM(15896) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(15896))))  severity failure;
	assert RAM(15897) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(15897))))  severity failure;
	assert RAM(15898) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(15898))))  severity failure;
	assert RAM(15899) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(15899))))  severity failure;
	assert RAM(15900) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(15900))))  severity failure;
	assert RAM(15901) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(15901))))  severity failure;
	assert RAM(15902) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(15902))))  severity failure;
	assert RAM(15903) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(15903))))  severity failure;
	assert RAM(15904) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(15904))))  severity failure;
	assert RAM(15905) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(15905))))  severity failure;
	assert RAM(15906) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(15906))))  severity failure;
	assert RAM(15907) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(15907))))  severity failure;
	assert RAM(15908) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(15908))))  severity failure;
	assert RAM(15909) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(15909))))  severity failure;
	assert RAM(15910) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(15910))))  severity failure;
	assert RAM(15911) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(15911))))  severity failure;
	assert RAM(15912) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(15912))))  severity failure;
	assert RAM(15913) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15913))))  severity failure;
	assert RAM(15914) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(15914))))  severity failure;
	assert RAM(15915) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(15915))))  severity failure;
	assert RAM(15916) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(15916))))  severity failure;
	assert RAM(15917) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(15917))))  severity failure;
	assert RAM(15918) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(15918))))  severity failure;
	assert RAM(15919) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(15919))))  severity failure;
	assert RAM(15920) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(15920))))  severity failure;
	assert RAM(15921) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(15921))))  severity failure;
	assert RAM(15922) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(15922))))  severity failure;
	assert RAM(15923) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(15923))))  severity failure;
	assert RAM(15924) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(15924))))  severity failure;
	assert RAM(15925) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(15925))))  severity failure;
	assert RAM(15926) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(15926))))  severity failure;
	assert RAM(15927) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(15927))))  severity failure;
	assert RAM(15928) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(15928))))  severity failure;
	assert RAM(15929) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(15929))))  severity failure;
	assert RAM(15930) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(15930))))  severity failure;
	assert RAM(15931) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(15931))))  severity failure;
	assert RAM(15932) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(15932))))  severity failure;
	assert RAM(15933) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(15933))))  severity failure;
	assert RAM(15934) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(15934))))  severity failure;
	assert RAM(15935) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(15935))))  severity failure;
	assert RAM(15936) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(15936))))  severity failure;
	assert RAM(15937) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(15937))))  severity failure;
	assert RAM(15938) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(15938))))  severity failure;
	assert RAM(15939) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(15939))))  severity failure;
	assert RAM(15940) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(15940))))  severity failure;
	assert RAM(15941) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(15941))))  severity failure;
	assert RAM(15942) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(15942))))  severity failure;
	assert RAM(15943) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(15943))))  severity failure;
	assert RAM(15944) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(15944))))  severity failure;
	assert RAM(15945) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(15945))))  severity failure;
	assert RAM(15946) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(15946))))  severity failure;
	assert RAM(15947) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(15947))))  severity failure;
	assert RAM(15948) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(15948))))  severity failure;
	assert RAM(15949) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(15949))))  severity failure;
	assert RAM(15950) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(15950))))  severity failure;
	assert RAM(15951) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(15951))))  severity failure;
	assert RAM(15952) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(15952))))  severity failure;
	assert RAM(15953) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(15953))))  severity failure;
	assert RAM(15954) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(15954))))  severity failure;
	assert RAM(15955) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(15955))))  severity failure;
	assert RAM(15956) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(15956))))  severity failure;
	assert RAM(15957) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(15957))))  severity failure;
	assert RAM(15958) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(15958))))  severity failure;
	assert RAM(15959) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(15959))))  severity failure;
	assert RAM(15960) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(15960))))  severity failure;
	assert RAM(15961) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(15961))))  severity failure;
	assert RAM(15962) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(15962))))  severity failure;
	assert RAM(15963) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(15963))))  severity failure;
	assert RAM(15964) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(15964))))  severity failure;
	assert RAM(15965) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(15965))))  severity failure;
	assert RAM(15966) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(15966))))  severity failure;
	assert RAM(15967) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(15967))))  severity failure;
	assert RAM(15968) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(15968))))  severity failure;
	assert RAM(15969) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(15969))))  severity failure;
	assert RAM(15970) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(15970))))  severity failure;
	assert RAM(15971) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(15971))))  severity failure;
	assert RAM(15972) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(15972))))  severity failure;
	assert RAM(15973) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(15973))))  severity failure;
	assert RAM(15974) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(15974))))  severity failure;
	assert RAM(15975) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(15975))))  severity failure;
	assert RAM(15976) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(15976))))  severity failure;
	assert RAM(15977) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(15977))))  severity failure;
	assert RAM(15978) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(15978))))  severity failure;
	assert RAM(15979) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(15979))))  severity failure;
	assert RAM(15980) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(15980))))  severity failure;
	assert RAM(15981) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(15981))))  severity failure;
	assert RAM(15982) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(15982))))  severity failure;
	assert RAM(15983) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(15983))))  severity failure;
	assert RAM(15984) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(15984))))  severity failure;
	assert RAM(15985) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(15985))))  severity failure;
	assert RAM(15986) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(15986))))  severity failure;
	assert RAM(15987) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(15987))))  severity failure;
	assert RAM(15988) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(15988))))  severity failure;
	assert RAM(15989) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(15989))))  severity failure;
	assert RAM(15990) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(15990))))  severity failure;
	assert RAM(15991) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(15991))))  severity failure;
	assert RAM(15992) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(15992))))  severity failure;
	assert RAM(15993) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(15993))))  severity failure;
	assert RAM(15994) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(15994))))  severity failure;
	assert RAM(15995) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(15995))))  severity failure;
	assert RAM(15996) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(15996))))  severity failure;
	assert RAM(15997) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(15997))))  severity failure;
	assert RAM(15998) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(15998))))  severity failure;
	assert RAM(15999) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(15999))))  severity failure;
	assert RAM(16000) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(16000))))  severity failure;
	assert RAM(16001) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(16001))))  severity failure;
	assert RAM(16002) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(16002))))  severity failure;
	assert RAM(16003) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16003))))  severity failure;
	assert RAM(16004) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(16004))))  severity failure;
	assert RAM(16005) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(16005))))  severity failure;
	assert RAM(16006) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(16006))))  severity failure;
	assert RAM(16007) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(16007))))  severity failure;
	assert RAM(16008) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(16008))))  severity failure;
	assert RAM(16009) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(16009))))  severity failure;
	assert RAM(16010) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(16010))))  severity failure;
	assert RAM(16011) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(16011))))  severity failure;
	assert RAM(16012) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(16012))))  severity failure;
	assert RAM(16013) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(16013))))  severity failure;
	assert RAM(16014) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16014))))  severity failure;
	assert RAM(16015) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(16015))))  severity failure;
	assert RAM(16016) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(16016))))  severity failure;
	assert RAM(16017) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(16017))))  severity failure;
	assert RAM(16018) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(16018))))  severity failure;
	assert RAM(16019) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(16019))))  severity failure;
	assert RAM(16020) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(16020))))  severity failure;
	assert RAM(16021) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(16021))))  severity failure;
	assert RAM(16022) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(16022))))  severity failure;
	assert RAM(16023) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16023))))  severity failure;
	assert RAM(16024) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(16024))))  severity failure;
	assert RAM(16025) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(16025))))  severity failure;
	assert RAM(16026) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(16026))))  severity failure;
	assert RAM(16027) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(16027))))  severity failure;
	assert RAM(16028) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(16028))))  severity failure;
	assert RAM(16029) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(16029))))  severity failure;
	assert RAM(16030) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(16030))))  severity failure;
	assert RAM(16031) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(16031))))  severity failure;
	assert RAM(16032) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(16032))))  severity failure;
	assert RAM(16033) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(16033))))  severity failure;
	assert RAM(16034) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(16034))))  severity failure;
	assert RAM(16035) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(16035))))  severity failure;
	assert RAM(16036) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(16036))))  severity failure;
	assert RAM(16037) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16037))))  severity failure;
	assert RAM(16038) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(16038))))  severity failure;
	assert RAM(16039) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(16039))))  severity failure;
	assert RAM(16040) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(16040))))  severity failure;
	assert RAM(16041) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(16041))))  severity failure;
	assert RAM(16042) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(16042))))  severity failure;
	assert RAM(16043) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(16043))))  severity failure;
	assert RAM(16044) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(16044))))  severity failure;
	assert RAM(16045) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(16045))))  severity failure;
	assert RAM(16046) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(16046))))  severity failure;
	assert RAM(16047) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(16047))))  severity failure;
	assert RAM(16048) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(16048))))  severity failure;
	assert RAM(16049) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(16049))))  severity failure;
	assert RAM(16050) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(16050))))  severity failure;
	assert RAM(16051) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(16051))))  severity failure;
	assert RAM(16052) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(16052))))  severity failure;
	assert RAM(16053) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(16053))))  severity failure;
	assert RAM(16054) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(16054))))  severity failure;
	assert RAM(16055) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(16055))))  severity failure;
	assert RAM(16056) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(16056))))  severity failure;
	assert RAM(16057) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(16057))))  severity failure;
	assert RAM(16058) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(16058))))  severity failure;
	assert RAM(16059) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(16059))))  severity failure;
	assert RAM(16060) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(16060))))  severity failure;
	assert RAM(16061) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16061))))  severity failure;
	assert RAM(16062) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(16062))))  severity failure;
	assert RAM(16063) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(16063))))  severity failure;
	assert RAM(16064) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(16064))))  severity failure;
	assert RAM(16065) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16065))))  severity failure;
	assert RAM(16066) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(16066))))  severity failure;
	assert RAM(16067) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(16067))))  severity failure;
	assert RAM(16068) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(16068))))  severity failure;
	assert RAM(16069) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16069))))  severity failure;
	assert RAM(16070) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16070))))  severity failure;
	assert RAM(16071) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16071))))  severity failure;
	assert RAM(16072) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(16072))))  severity failure;
	assert RAM(16073) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(16073))))  severity failure;
	assert RAM(16074) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(16074))))  severity failure;
	assert RAM(16075) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(16075))))  severity failure;
	assert RAM(16076) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(16076))))  severity failure;
	assert RAM(16077) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(16077))))  severity failure;
	assert RAM(16078) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(16078))))  severity failure;
	assert RAM(16079) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(16079))))  severity failure;
	assert RAM(16080) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(16080))))  severity failure;
	assert RAM(16081) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(16081))))  severity failure;
	assert RAM(16082) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(16082))))  severity failure;
	assert RAM(16083) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16083))))  severity failure;
	assert RAM(16084) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(16084))))  severity failure;
	assert RAM(16085) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16085))))  severity failure;
	assert RAM(16086) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(16086))))  severity failure;
	assert RAM(16087) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16087))))  severity failure;
	assert RAM(16088) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(16088))))  severity failure;
	assert RAM(16089) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(16089))))  severity failure;
	assert RAM(16090) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(16090))))  severity failure;
	assert RAM(16091) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16091))))  severity failure;
	assert RAM(16092) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(16092))))  severity failure;
	assert RAM(16093) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(16093))))  severity failure;
	assert RAM(16094) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(16094))))  severity failure;
	assert RAM(16095) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(16095))))  severity failure;
	assert RAM(16096) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(16096))))  severity failure;
	assert RAM(16097) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16097))))  severity failure;
	assert RAM(16098) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(16098))))  severity failure;
	assert RAM(16099) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(16099))))  severity failure;
	assert RAM(16100) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(16100))))  severity failure;
	assert RAM(16101) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(16101))))  severity failure;
	assert RAM(16102) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(16102))))  severity failure;
	assert RAM(16103) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(16103))))  severity failure;
	assert RAM(16104) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(16104))))  severity failure;
	assert RAM(16105) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(16105))))  severity failure;
	assert RAM(16106) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(16106))))  severity failure;
	assert RAM(16107) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(16107))))  severity failure;
	assert RAM(16108) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(16108))))  severity failure;
	assert RAM(16109) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(16109))))  severity failure;
	assert RAM(16110) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(16110))))  severity failure;
	assert RAM(16111) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16111))))  severity failure;
	assert RAM(16112) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(16112))))  severity failure;
	assert RAM(16113) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(16113))))  severity failure;
	assert RAM(16114) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(16114))))  severity failure;
	assert RAM(16115) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(16115))))  severity failure;
	assert RAM(16116) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(16116))))  severity failure;
	assert RAM(16117) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(16117))))  severity failure;
	assert RAM(16118) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(16118))))  severity failure;
	assert RAM(16119) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(16119))))  severity failure;
	assert RAM(16120) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(16120))))  severity failure;
	assert RAM(16121) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(16121))))  severity failure;
	assert RAM(16122) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(16122))))  severity failure;
	assert RAM(16123) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16123))))  severity failure;
	assert RAM(16124) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(16124))))  severity failure;
	assert RAM(16125) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16125))))  severity failure;
	assert RAM(16126) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16126))))  severity failure;
	assert RAM(16127) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(16127))))  severity failure;
	assert RAM(16128) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(16128))))  severity failure;
	assert RAM(16129) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(16129))))  severity failure;
	assert RAM(16130) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16130))))  severity failure;
	assert RAM(16131) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16131))))  severity failure;
	assert RAM(16132) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(16132))))  severity failure;
	assert RAM(16133) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16133))))  severity failure;
	assert RAM(16134) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(16134))))  severity failure;
	assert RAM(16135) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16135))))  severity failure;
	assert RAM(16136) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(16136))))  severity failure;
	assert RAM(16137) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(16137))))  severity failure;
	assert RAM(16138) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(16138))))  severity failure;
	assert RAM(16139) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(16139))))  severity failure;
	assert RAM(16140) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(16140))))  severity failure;
	assert RAM(16141) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(16141))))  severity failure;
	assert RAM(16142) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(16142))))  severity failure;
	assert RAM(16143) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(16143))))  severity failure;
	assert RAM(16144) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(16144))))  severity failure;
	assert RAM(16145) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16145))))  severity failure;
	assert RAM(16146) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(16146))))  severity failure;
	assert RAM(16147) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(16147))))  severity failure;
	assert RAM(16148) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(16148))))  severity failure;
	assert RAM(16149) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16149))))  severity failure;
	assert RAM(16150) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(16150))))  severity failure;
	assert RAM(16151) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(16151))))  severity failure;
	assert RAM(16152) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(16152))))  severity failure;
	assert RAM(16153) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(16153))))  severity failure;
	assert RAM(16154) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(16154))))  severity failure;
	assert RAM(16155) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(16155))))  severity failure;
	assert RAM(16156) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(16156))))  severity failure;
	assert RAM(16157) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(16157))))  severity failure;
	assert RAM(16158) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(16158))))  severity failure;
	assert RAM(16159) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(16159))))  severity failure;
	assert RAM(16160) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(16160))))  severity failure;
	assert RAM(16161) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(16161))))  severity failure;
	assert RAM(16162) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(16162))))  severity failure;
	assert RAM(16163) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(16163))))  severity failure;
	assert RAM(16164) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(16164))))  severity failure;
	assert RAM(16165) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(16165))))  severity failure;
	assert RAM(16166) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(16166))))  severity failure;
	assert RAM(16167) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(16167))))  severity failure;
	assert RAM(16168) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(16168))))  severity failure;
	assert RAM(16169) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(16169))))  severity failure;
	assert RAM(16170) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(16170))))  severity failure;
	assert RAM(16171) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(16171))))  severity failure;
	assert RAM(16172) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(16172))))  severity failure;
	assert RAM(16173) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16173))))  severity failure;
	assert RAM(16174) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(16174))))  severity failure;
	assert RAM(16175) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(16175))))  severity failure;
	assert RAM(16176) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(16176))))  severity failure;
	assert RAM(16177) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(16177))))  severity failure;
	assert RAM(16178) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(16178))))  severity failure;
	assert RAM(16179) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(16179))))  severity failure;
	assert RAM(16180) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(16180))))  severity failure;
	assert RAM(16181) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(16181))))  severity failure;
	assert RAM(16182) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(16182))))  severity failure;
	assert RAM(16183) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(16183))))  severity failure;
	assert RAM(16184) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(16184))))  severity failure;
	assert RAM(16185) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(16185))))  severity failure;
	assert RAM(16186) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(16186))))  severity failure;
	assert RAM(16187) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(16187))))  severity failure;
	assert RAM(16188) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(16188))))  severity failure;
	assert RAM(16189) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(16189))))  severity failure;
	assert RAM(16190) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(16190))))  severity failure;
	assert RAM(16191) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(16191))))  severity failure;
	assert RAM(16192) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16192))))  severity failure;
	assert RAM(16193) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(16193))))  severity failure;
	assert RAM(16194) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(16194))))  severity failure;
	assert RAM(16195) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(16195))))  severity failure;
	assert RAM(16196) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(16196))))  severity failure;
	assert RAM(16197) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(16197))))  severity failure;
	assert RAM(16198) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(16198))))  severity failure;
	assert RAM(16199) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(16199))))  severity failure;
	assert RAM(16200) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16200))))  severity failure;
	assert RAM(16201) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(16201))))  severity failure;
	assert RAM(16202) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16202))))  severity failure;
	assert RAM(16203) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(16203))))  severity failure;
	assert RAM(16204) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(16204))))  severity failure;
	assert RAM(16205) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(16205))))  severity failure;
	assert RAM(16206) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(16206))))  severity failure;
	assert RAM(16207) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(16207))))  severity failure;
	assert RAM(16208) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16208))))  severity failure;
	assert RAM(16209) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16209))))  severity failure;
	assert RAM(16210) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(16210))))  severity failure;
	assert RAM(16211) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(16211))))  severity failure;
	assert RAM(16212) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16212))))  severity failure;
	assert RAM(16213) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(16213))))  severity failure;
	assert RAM(16214) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16214))))  severity failure;
	assert RAM(16215) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(16215))))  severity failure;
	assert RAM(16216) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(16216))))  severity failure;
	assert RAM(16217) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(16217))))  severity failure;
	assert RAM(16218) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(16218))))  severity failure;
	assert RAM(16219) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(16219))))  severity failure;
	assert RAM(16220) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(16220))))  severity failure;
	assert RAM(16221) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(16221))))  severity failure;
	assert RAM(16222) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(16222))))  severity failure;
	assert RAM(16223) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(16223))))  severity failure;
	assert RAM(16224) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(16224))))  severity failure;
	assert RAM(16225) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(16225))))  severity failure;
	assert RAM(16226) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(16226))))  severity failure;
	assert RAM(16227) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16227))))  severity failure;
	assert RAM(16228) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(16228))))  severity failure;
	assert RAM(16229) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(16229))))  severity failure;
	assert RAM(16230) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(16230))))  severity failure;
	assert RAM(16231) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(16231))))  severity failure;
	assert RAM(16232) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(16232))))  severity failure;
	assert RAM(16233) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(16233))))  severity failure;
	assert RAM(16234) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(16234))))  severity failure;
	assert RAM(16235) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(16235))))  severity failure;
	assert RAM(16236) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(16236))))  severity failure;
	assert RAM(16237) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(16237))))  severity failure;
	assert RAM(16238) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16238))))  severity failure;
	assert RAM(16239) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(16239))))  severity failure;
	assert RAM(16240) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(16240))))  severity failure;
	assert RAM(16241) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(16241))))  severity failure;
	assert RAM(16242) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(16242))))  severity failure;
	assert RAM(16243) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(16243))))  severity failure;
	assert RAM(16244) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(16244))))  severity failure;
	assert RAM(16245) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(16245))))  severity failure;
	assert RAM(16246) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16246))))  severity failure;
	assert RAM(16247) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(16247))))  severity failure;
	assert RAM(16248) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(16248))))  severity failure;
	assert RAM(16249) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(16249))))  severity failure;
	assert RAM(16250) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16250))))  severity failure;
	assert RAM(16251) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(16251))))  severity failure;
	assert RAM(16252) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(16252))))  severity failure;
	assert RAM(16253) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(16253))))  severity failure;
	assert RAM(16254) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(16254))))  severity failure;
	assert RAM(16255) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(16255))))  severity failure;
	assert RAM(16256) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(16256))))  severity failure;
	assert RAM(16257) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(16257))))  severity failure;
	assert RAM(16258) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(16258))))  severity failure;
	assert RAM(16259) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(16259))))  severity failure;
	assert RAM(16260) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(16260))))  severity failure;
	assert RAM(16261) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(16261))))  severity failure;
	assert RAM(16262) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(16262))))  severity failure;
	assert RAM(16263) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(16263))))  severity failure;
	assert RAM(16264) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(16264))))  severity failure;
	assert RAM(16265) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16265))))  severity failure;
	assert RAM(16266) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(16266))))  severity failure;
	assert RAM(16267) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(16267))))  severity failure;
	assert RAM(16268) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16268))))  severity failure;
	assert RAM(16269) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16269))))  severity failure;
	assert RAM(16270) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(16270))))  severity failure;
	assert RAM(16271) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(16271))))  severity failure;
	assert RAM(16272) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(16272))))  severity failure;
	assert RAM(16273) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(16273))))  severity failure;
	assert RAM(16274) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(16274))))  severity failure;
	assert RAM(16275) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(16275))))  severity failure;
	assert RAM(16276) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(16276))))  severity failure;
	assert RAM(16277) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(16277))))  severity failure;
	assert RAM(16278) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16278))))  severity failure;
	assert RAM(16279) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(16279))))  severity failure;
	assert RAM(16280) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(16280))))  severity failure;
	assert RAM(16281) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(16281))))  severity failure;
	assert RAM(16282) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(16282))))  severity failure;
	assert RAM(16283) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(16283))))  severity failure;
	assert RAM(16284) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(16284))))  severity failure;
	assert RAM(16285) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16285))))  severity failure;
	assert RAM(16286) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(16286))))  severity failure;
	assert RAM(16287) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(16287))))  severity failure;
	assert RAM(16288) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(16288))))  severity failure;
	assert RAM(16289) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(16289))))  severity failure;
	assert RAM(16290) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16290))))  severity failure;
	assert RAM(16291) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(16291))))  severity failure;
	assert RAM(16292) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(16292))))  severity failure;
	assert RAM(16293) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(16293))))  severity failure;
	assert RAM(16294) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(16294))))  severity failure;
	assert RAM(16295) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(16295))))  severity failure;
	assert RAM(16296) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(16296))))  severity failure;
	assert RAM(16297) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(16297))))  severity failure;
	assert RAM(16298) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(16298))))  severity failure;
	assert RAM(16299) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(16299))))  severity failure;
	assert RAM(16300) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(16300))))  severity failure;
	assert RAM(16301) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(16301))))  severity failure;
	assert RAM(16302) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(16302))))  severity failure;
	assert RAM(16303) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(16303))))  severity failure;
	assert RAM(16304) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(16304))))  severity failure;
	assert RAM(16305) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(16305))))  severity failure;
	assert RAM(16306) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(16306))))  severity failure;
	assert RAM(16307) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(16307))))  severity failure;
	assert RAM(16308) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16308))))  severity failure;
	assert RAM(16309) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(16309))))  severity failure;
	assert RAM(16310) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(16310))))  severity failure;
	assert RAM(16311) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(16311))))  severity failure;
	assert RAM(16312) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(16312))))  severity failure;
	assert RAM(16313) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(16313))))  severity failure;
	assert RAM(16314) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(16314))))  severity failure;
	assert RAM(16315) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(16315))))  severity failure;
	assert RAM(16316) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(16316))))  severity failure;
	assert RAM(16317) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(16317))))  severity failure;
	assert RAM(16318) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16318))))  severity failure;
	assert RAM(16319) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(16319))))  severity failure;
	assert RAM(16320) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(16320))))  severity failure;
	assert RAM(16321) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16321))))  severity failure;
	assert RAM(16322) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(16322))))  severity failure;
	assert RAM(16323) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(16323))))  severity failure;
	assert RAM(16324) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(16324))))  severity failure;
	assert RAM(16325) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(16325))))  severity failure;
	assert RAM(16326) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(16326))))  severity failure;
	assert RAM(16327) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(16327))))  severity failure;
	assert RAM(16328) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(16328))))  severity failure;
	assert RAM(16329) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(16329))))  severity failure;
	assert RAM(16330) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16330))))  severity failure;
	assert RAM(16331) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(16331))))  severity failure;
	assert RAM(16332) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(16332))))  severity failure;
	assert RAM(16333) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(16333))))  severity failure;
	assert RAM(16334) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(16334))))  severity failure;
	assert RAM(16335) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(16335))))  severity failure;
	assert RAM(16336) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16336))))  severity failure;
	assert RAM(16337) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(16337))))  severity failure;
	assert RAM(16338) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16338))))  severity failure;
	assert RAM(16339) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(16339))))  severity failure;
	assert RAM(16340) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(16340))))  severity failure;
	assert RAM(16341) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(16341))))  severity failure;
	assert RAM(16342) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(16342))))  severity failure;
	assert RAM(16343) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(16343))))  severity failure;
	assert RAM(16344) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(16344))))  severity failure;
	assert RAM(16345) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(16345))))  severity failure;
	assert RAM(16346) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(16346))))  severity failure;
	assert RAM(16347) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16347))))  severity failure;
	assert RAM(16348) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(16348))))  severity failure;
	assert RAM(16349) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(16349))))  severity failure;
	assert RAM(16350) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(16350))))  severity failure;
	assert RAM(16351) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(16351))))  severity failure;
	assert RAM(16352) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(16352))))  severity failure;
	assert RAM(16353) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(16353))))  severity failure;
	assert RAM(16354) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(16354))))  severity failure;
	assert RAM(16355) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(16355))))  severity failure;
	assert RAM(16356) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16356))))  severity failure;
	assert RAM(16357) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(16357))))  severity failure;
	assert RAM(16358) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(16358))))  severity failure;
	assert RAM(16359) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(16359))))  severity failure;
	assert RAM(16360) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(16360))))  severity failure;
	assert RAM(16361) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(16361))))  severity failure;
	assert RAM(16362) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(16362))))  severity failure;
	assert RAM(16363) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(16363))))  severity failure;
	assert RAM(16364) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16364))))  severity failure;
	assert RAM(16365) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(16365))))  severity failure;
	assert RAM(16366) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(16366))))  severity failure;
	assert RAM(16367) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(16367))))  severity failure;
	assert RAM(16368) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16368))))  severity failure;
	assert RAM(16369) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16369))))  severity failure;
	assert RAM(16370) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(16370))))  severity failure;
	assert RAM(16371) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(16371))))  severity failure;
	assert RAM(16372) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(16372))))  severity failure;
	assert RAM(16373) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(16373))))  severity failure;
	assert RAM(16374) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(16374))))  severity failure;
	assert RAM(16375) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(16375))))  severity failure;
	assert RAM(16376) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(16376))))  severity failure;
	assert RAM(16377) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(16377))))  severity failure;
	assert RAM(16378) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(16378))))  severity failure;
	assert RAM(16379) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(16379))))  severity failure;
	assert RAM(16380) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(16380))))  severity failure;
	assert RAM(16381) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(16381))))  severity failure;
	assert RAM(16382) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(16382))))  severity failure;
	assert RAM(16383) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(16383))))  severity failure;
	assert RAM(16384) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(16384))))  severity failure;
	assert RAM(16385) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(16385))))  severity failure;
	assert RAM(16386) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(16386))))  severity failure;
	assert RAM(16387) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16387))))  severity failure;
	assert RAM(16388) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(16388))))  severity failure;
	assert RAM(16389) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(16389))))  severity failure;
	assert RAM(16390) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(16390))))  severity failure;
	assert RAM(16391) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(16391))))  severity failure;
	assert RAM(16392) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(16392))))  severity failure;
	assert RAM(16393) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(16393))))  severity failure;
	assert RAM(16394) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(16394))))  severity failure;
	assert RAM(16395) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(16395))))  severity failure;
	assert RAM(16396) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(16396))))  severity failure;
	assert RAM(16397) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(16397))))  severity failure;
	assert RAM(16398) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(16398))))  severity failure;
	assert RAM(16399) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(16399))))  severity failure;
	assert RAM(16400) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(16400))))  severity failure;
	assert RAM(16401) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(16401))))  severity failure;
	assert RAM(16402) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(16402))))  severity failure;
	assert RAM(16403) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(16403))))  severity failure;
	assert RAM(16404) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(16404))))  severity failure;
	assert RAM(16405) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(16405))))  severity failure;
	assert RAM(16406) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(16406))))  severity failure;
	assert RAM(16407) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(16407))))  severity failure;
	assert RAM(16408) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(16408))))  severity failure;
	assert RAM(16409) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16409))))  severity failure;
	assert RAM(16410) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(16410))))  severity failure;
	assert RAM(16411) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16411))))  severity failure;
	assert RAM(16412) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(16412))))  severity failure;
	assert RAM(16413) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(16413))))  severity failure;
	assert RAM(16414) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(16414))))  severity failure;
	assert RAM(16415) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(16415))))  severity failure;
	assert RAM(16416) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(16416))))  severity failure;
	assert RAM(16417) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(16417))))  severity failure;
	assert RAM(16418) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(16418))))  severity failure;
	assert RAM(16419) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16419))))  severity failure;
	assert RAM(16420) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(16420))))  severity failure;
	assert RAM(16421) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(16421))))  severity failure;
	assert RAM(16422) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(16422))))  severity failure;
	assert RAM(16423) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(16423))))  severity failure;
	assert RAM(16424) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(16424))))  severity failure;
	assert RAM(16425) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(16425))))  severity failure;
	assert RAM(16426) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(16426))))  severity failure;
	assert RAM(16427) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(16427))))  severity failure;
	assert RAM(16428) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(16428))))  severity failure;
	assert RAM(16429) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(16429))))  severity failure;
	assert RAM(16430) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(16430))))  severity failure;
	assert RAM(16431) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(16431))))  severity failure;
	assert RAM(16432) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(16432))))  severity failure;
	assert RAM(16433) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(16433))))  severity failure;
	assert RAM(16434) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(16434))))  severity failure;
	assert RAM(16435) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(16435))))  severity failure;
	assert RAM(16436) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(16436))))  severity failure;
	assert RAM(16437) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(16437))))  severity failure;
	assert RAM(16438) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(16438))))  severity failure;
	assert RAM(16439) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(16439))))  severity failure;
	assert RAM(16440) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(16440))))  severity failure;
	assert RAM(16441) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(16441))))  severity failure;
	assert RAM(16442) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(16442))))  severity failure;
	assert RAM(16443) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(16443))))  severity failure;
	assert RAM(16444) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(16444))))  severity failure;
	assert RAM(16445) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(16445))))  severity failure;
	assert RAM(16446) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(16446))))  severity failure;
	assert RAM(16447) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(16447))))  severity failure;
	assert RAM(16448) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(16448))))  severity failure;
	assert RAM(16449) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16449))))  severity failure;
	assert RAM(16450) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(16450))))  severity failure;
	assert RAM(16451) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(16451))))  severity failure;
	assert RAM(16452) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(16452))))  severity failure;
	assert RAM(16453) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(16453))))  severity failure;
	assert RAM(16454) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(16454))))  severity failure;
	assert RAM(16455) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(16455))))  severity failure;
	assert RAM(16456) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(16456))))  severity failure;
	assert RAM(16457) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(16457))))  severity failure;
	assert RAM(16458) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(16458))))  severity failure;
	assert RAM(16459) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(16459))))  severity failure;
	assert RAM(16460) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(16460))))  severity failure;
	assert RAM(16461) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(16461))))  severity failure;
	assert RAM(16462) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(16462))))  severity failure;
	assert RAM(16463) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16463))))  severity failure;
	assert RAM(16464) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(16464))))  severity failure;
	assert RAM(16465) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(16465))))  severity failure;
	assert RAM(16466) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(16466))))  severity failure;
	assert RAM(16467) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(16467))))  severity failure;
	assert RAM(16468) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(16468))))  severity failure;
	assert RAM(16469) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(16469))))  severity failure;
	assert RAM(16470) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(16470))))  severity failure;
	assert RAM(16471) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(16471))))  severity failure;
	assert RAM(16472) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(16472))))  severity failure;
	assert RAM(16473) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(16473))))  severity failure;
	assert RAM(16474) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(16474))))  severity failure;
	assert RAM(16475) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(16475))))  severity failure;
	assert RAM(16476) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(16476))))  severity failure;
	assert RAM(16477) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(16477))))  severity failure;
	assert RAM(16478) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(16478))))  severity failure;
	assert RAM(16479) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(16479))))  severity failure;
	assert RAM(16480) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(16480))))  severity failure;
	assert RAM(16481) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(16481))))  severity failure;
	assert RAM(16482) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(16482))))  severity failure;
	assert RAM(16483) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(16483))))  severity failure;
	assert RAM(16484) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(16484))))  severity failure;
	assert RAM(16485) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(16485))))  severity failure;
	assert RAM(16486) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(16486))))  severity failure;
	assert RAM(16487) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(16487))))  severity failure;
	assert RAM(16488) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16488))))  severity failure;
	assert RAM(16489) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(16489))))  severity failure;
	assert RAM(16490) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(16490))))  severity failure;
	assert RAM(16491) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(16491))))  severity failure;
	assert RAM(16492) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(16492))))  severity failure;
	assert RAM(16493) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(16493))))  severity failure;
	assert RAM(16494) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(16494))))  severity failure;
	assert RAM(16495) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(16495))))  severity failure;
	assert RAM(16496) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(16496))))  severity failure;
	assert RAM(16497) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16497))))  severity failure;
	assert RAM(16498) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16498))))  severity failure;
	assert RAM(16499) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(16499))))  severity failure;
	assert RAM(16500) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16500))))  severity failure;
	assert RAM(16501) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(16501))))  severity failure;
	assert RAM(16502) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(16502))))  severity failure;
	assert RAM(16503) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(16503))))  severity failure;
	assert RAM(16504) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(16504))))  severity failure;
	assert RAM(16505) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(16505))))  severity failure;
	assert RAM(16506) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(16506))))  severity failure;
	assert RAM(16507) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(16507))))  severity failure;
	assert RAM(16508) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16508))))  severity failure;
	assert RAM(16509) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(16509))))  severity failure;
	assert RAM(16510) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(16510))))  severity failure;
	assert RAM(16511) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(16511))))  severity failure;
	assert RAM(16512) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16512))))  severity failure;
	assert RAM(16513) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(16513))))  severity failure;
	assert RAM(16514) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(16514))))  severity failure;
	assert RAM(16515) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(16515))))  severity failure;
	assert RAM(16516) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(16516))))  severity failure;
	assert RAM(16517) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(16517))))  severity failure;
	assert RAM(16518) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(16518))))  severity failure;
	assert RAM(16519) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(16519))))  severity failure;
	assert RAM(16520) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(16520))))  severity failure;
	assert RAM(16521) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(16521))))  severity failure;
	assert RAM(16522) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(16522))))  severity failure;
	assert RAM(16523) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16523))))  severity failure;
	assert RAM(16524) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(16524))))  severity failure;
	assert RAM(16525) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(16525))))  severity failure;
	assert RAM(16526) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(16526))))  severity failure;
	assert RAM(16527) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(16527))))  severity failure;
	assert RAM(16528) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16528))))  severity failure;
	assert RAM(16529) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(16529))))  severity failure;
	assert RAM(16530) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(16530))))  severity failure;
	assert RAM(16531) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(16531))))  severity failure;
	assert RAM(16532) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(16532))))  severity failure;
	assert RAM(16533) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(16533))))  severity failure;
	assert RAM(16534) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(16534))))  severity failure;
	assert RAM(16535) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(16535))))  severity failure;
	assert RAM(16536) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(16536))))  severity failure;
	assert RAM(16537) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(16537))))  severity failure;
	assert RAM(16538) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(16538))))  severity failure;
	assert RAM(16539) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(16539))))  severity failure;
	assert RAM(16540) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(16540))))  severity failure;
	assert RAM(16541) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(16541))))  severity failure;
	assert RAM(16542) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16542))))  severity failure;
	assert RAM(16543) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(16543))))  severity failure;
	assert RAM(16544) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(16544))))  severity failure;
	assert RAM(16545) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(16545))))  severity failure;
	assert RAM(16546) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(16546))))  severity failure;
	assert RAM(16547) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(16547))))  severity failure;
	assert RAM(16548) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(16548))))  severity failure;
	assert RAM(16549) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(16549))))  severity failure;
	assert RAM(16550) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(16550))))  severity failure;
	assert RAM(16551) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16551))))  severity failure;
	assert RAM(16552) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16552))))  severity failure;
	assert RAM(16553) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16553))))  severity failure;
	assert RAM(16554) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16554))))  severity failure;
	assert RAM(16555) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(16555))))  severity failure;
	assert RAM(16556) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(16556))))  severity failure;
	assert RAM(16557) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(16557))))  severity failure;
	assert RAM(16558) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(16558))))  severity failure;
	assert RAM(16559) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(16559))))  severity failure;
	assert RAM(16560) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(16560))))  severity failure;
	assert RAM(16561) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(16561))))  severity failure;
	assert RAM(16562) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16562))))  severity failure;
	assert RAM(16563) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(16563))))  severity failure;
	assert RAM(16564) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(16564))))  severity failure;
	assert RAM(16565) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(16565))))  severity failure;
	assert RAM(16566) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16566))))  severity failure;
	assert RAM(16567) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(16567))))  severity failure;
	assert RAM(16568) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(16568))))  severity failure;
	assert RAM(16569) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(16569))))  severity failure;
	assert RAM(16570) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(16570))))  severity failure;
	assert RAM(16571) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(16571))))  severity failure;
	assert RAM(16572) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(16572))))  severity failure;
	assert RAM(16573) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(16573))))  severity failure;
	assert RAM(16574) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(16574))))  severity failure;
	assert RAM(16575) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(16575))))  severity failure;
	assert RAM(16576) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(16576))))  severity failure;
	assert RAM(16577) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(16577))))  severity failure;
	assert RAM(16578) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(16578))))  severity failure;
	assert RAM(16579) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(16579))))  severity failure;
	assert RAM(16580) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(16580))))  severity failure;
	assert RAM(16581) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(16581))))  severity failure;
	assert RAM(16582) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(16582))))  severity failure;
	assert RAM(16583) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(16583))))  severity failure;
	assert RAM(16584) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(16584))))  severity failure;
	assert RAM(16585) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(16585))))  severity failure;
	assert RAM(16586) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(16586))))  severity failure;
	assert RAM(16587) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(16587))))  severity failure;
	assert RAM(16588) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(16588))))  severity failure;
	assert RAM(16589) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(16589))))  severity failure;
	assert RAM(16590) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(16590))))  severity failure;
	assert RAM(16591) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(16591))))  severity failure;
	assert RAM(16592) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(16592))))  severity failure;
	assert RAM(16593) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(16593))))  severity failure;
	assert RAM(16594) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(16594))))  severity failure;
	assert RAM(16595) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(16595))))  severity failure;
	assert RAM(16596) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16596))))  severity failure;
	assert RAM(16597) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(16597))))  severity failure;
	assert RAM(16598) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(16598))))  severity failure;
	assert RAM(16599) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(16599))))  severity failure;
	assert RAM(16600) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(16600))))  severity failure;
	assert RAM(16601) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(16601))))  severity failure;
	assert RAM(16602) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(16602))))  severity failure;
	assert RAM(16603) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(16603))))  severity failure;
	assert RAM(16604) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(16604))))  severity failure;
	assert RAM(16605) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(16605))))  severity failure;
	assert RAM(16606) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16606))))  severity failure;
	assert RAM(16607) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(16607))))  severity failure;
	assert RAM(16608) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16608))))  severity failure;
	assert RAM(16609) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16609))))  severity failure;
	assert RAM(16610) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(16610))))  severity failure;
	assert RAM(16611) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(16611))))  severity failure;
	assert RAM(16612) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(16612))))  severity failure;
	assert RAM(16613) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16613))))  severity failure;
	assert RAM(16614) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(16614))))  severity failure;
	assert RAM(16615) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(16615))))  severity failure;
	assert RAM(16616) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(16616))))  severity failure;
	assert RAM(16617) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16617))))  severity failure;
	assert RAM(16618) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(16618))))  severity failure;
	assert RAM(16619) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(16619))))  severity failure;
	assert RAM(16620) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16620))))  severity failure;
	assert RAM(16621) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(16621))))  severity failure;
	assert RAM(16622) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(16622))))  severity failure;
	assert RAM(16623) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(16623))))  severity failure;
	assert RAM(16624) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(16624))))  severity failure;
	assert RAM(16625) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(16625))))  severity failure;
	assert RAM(16626) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(16626))))  severity failure;
	assert RAM(16627) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(16627))))  severity failure;
	assert RAM(16628) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(16628))))  severity failure;
	assert RAM(16629) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(16629))))  severity failure;
	assert RAM(16630) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16630))))  severity failure;
	assert RAM(16631) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(16631))))  severity failure;
	assert RAM(16632) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(16632))))  severity failure;
	assert RAM(16633) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(16633))))  severity failure;
	assert RAM(16634) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(16634))))  severity failure;
	assert RAM(16635) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(16635))))  severity failure;
	assert RAM(16636) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(16636))))  severity failure;
	assert RAM(16637) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(16637))))  severity failure;
	assert RAM(16638) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(16638))))  severity failure;
	assert RAM(16639) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(16639))))  severity failure;
	assert RAM(16640) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(16640))))  severity failure;
	assert RAM(16641) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(16641))))  severity failure;
	assert RAM(16642) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(16642))))  severity failure;
	assert RAM(16643) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(16643))))  severity failure;
	assert RAM(16644) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(16644))))  severity failure;
	assert RAM(16645) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(16645))))  severity failure;
	assert RAM(16646) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(16646))))  severity failure;
	assert RAM(16647) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(16647))))  severity failure;
	assert RAM(16648) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(16648))))  severity failure;
	assert RAM(16649) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(16649))))  severity failure;
	assert RAM(16650) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(16650))))  severity failure;
	assert RAM(16651) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(16651))))  severity failure;
	assert RAM(16652) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(16652))))  severity failure;
	assert RAM(16653) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(16653))))  severity failure;
	assert RAM(16654) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(16654))))  severity failure;
	assert RAM(16655) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(16655))))  severity failure;
	assert RAM(16656) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16656))))  severity failure;
	assert RAM(16657) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(16657))))  severity failure;
	assert RAM(16658) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(16658))))  severity failure;
	assert RAM(16659) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16659))))  severity failure;
	assert RAM(16660) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(16660))))  severity failure;
	assert RAM(16661) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(16661))))  severity failure;
	assert RAM(16662) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(16662))))  severity failure;
	assert RAM(16663) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(16663))))  severity failure;
	assert RAM(16664) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(16664))))  severity failure;
	assert RAM(16665) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(16665))))  severity failure;
	assert RAM(16666) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(16666))))  severity failure;
	assert RAM(16667) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(16667))))  severity failure;
	assert RAM(16668) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(16668))))  severity failure;
	assert RAM(16669) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(16669))))  severity failure;
	assert RAM(16670) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(16670))))  severity failure;
	assert RAM(16671) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16671))))  severity failure;
	assert RAM(16672) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(16672))))  severity failure;
	assert RAM(16673) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16673))))  severity failure;
	assert RAM(16674) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(16674))))  severity failure;
	assert RAM(16675) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(16675))))  severity failure;
	assert RAM(16676) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(16676))))  severity failure;
	assert RAM(16677) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(16677))))  severity failure;
	assert RAM(16678) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(16678))))  severity failure;
	assert RAM(16679) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(16679))))  severity failure;
	assert RAM(16680) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(16680))))  severity failure;
	assert RAM(16681) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(16681))))  severity failure;
	assert RAM(16682) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(16682))))  severity failure;
	assert RAM(16683) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(16683))))  severity failure;
	assert RAM(16684) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(16684))))  severity failure;
	assert RAM(16685) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(16685))))  severity failure;
	assert RAM(16686) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(16686))))  severity failure;
	assert RAM(16687) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(16687))))  severity failure;
	assert RAM(16688) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16688))))  severity failure;
	assert RAM(16689) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(16689))))  severity failure;
	assert RAM(16690) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(16690))))  severity failure;
	assert RAM(16691) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(16691))))  severity failure;
	assert RAM(16692) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(16692))))  severity failure;
	assert RAM(16693) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(16693))))  severity failure;
	assert RAM(16694) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(16694))))  severity failure;
	assert RAM(16695) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(16695))))  severity failure;
	assert RAM(16696) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(16696))))  severity failure;
	assert RAM(16697) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16697))))  severity failure;
	assert RAM(16698) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(16698))))  severity failure;
	assert RAM(16699) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(16699))))  severity failure;
	assert RAM(16700) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(16700))))  severity failure;
	assert RAM(16701) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(16701))))  severity failure;
	assert RAM(16702) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(16702))))  severity failure;
	assert RAM(16703) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(16703))))  severity failure;
	assert RAM(16704) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(16704))))  severity failure;
	assert RAM(16705) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16705))))  severity failure;
	assert RAM(16706) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(16706))))  severity failure;
	assert RAM(16707) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(16707))))  severity failure;
	assert RAM(16708) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(16708))))  severity failure;
	assert RAM(16709) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(16709))))  severity failure;
	assert RAM(16710) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(16710))))  severity failure;
	assert RAM(16711) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(16711))))  severity failure;
	assert RAM(16712) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(16712))))  severity failure;
	assert RAM(16713) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(16713))))  severity failure;
	assert RAM(16714) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(16714))))  severity failure;
	assert RAM(16715) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(16715))))  severity failure;
	assert RAM(16716) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(16716))))  severity failure;
	assert RAM(16717) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(16717))))  severity failure;
	assert RAM(16718) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(16718))))  severity failure;
	assert RAM(16719) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(16719))))  severity failure;
	assert RAM(16720) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(16720))))  severity failure;
	assert RAM(16721) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(16721))))  severity failure;
	assert RAM(16722) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(16722))))  severity failure;
	assert RAM(16723) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(16723))))  severity failure;
	assert RAM(16724) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(16724))))  severity failure;
	assert RAM(16725) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(16725))))  severity failure;
	assert RAM(16726) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(16726))))  severity failure;
	assert RAM(16727) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(16727))))  severity failure;
	assert RAM(16728) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(16728))))  severity failure;
	assert RAM(16729) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(16729))))  severity failure;
	assert RAM(16730) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(16730))))  severity failure;
	assert RAM(16731) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(16731))))  severity failure;
	assert RAM(16732) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(16732))))  severity failure;
	assert RAM(16733) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(16733))))  severity failure;
	assert RAM(16734) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16734))))  severity failure;
	assert RAM(16735) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(16735))))  severity failure;
	assert RAM(16736) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(16736))))  severity failure;
	assert RAM(16737) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(16737))))  severity failure;
	assert RAM(16738) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(16738))))  severity failure;
	assert RAM(16739) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(16739))))  severity failure;
	assert RAM(16740) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(16740))))  severity failure;
	assert RAM(16741) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(16741))))  severity failure;
	assert RAM(16742) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(16742))))  severity failure;
	assert RAM(16743) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(16743))))  severity failure;
	assert RAM(16744) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(16744))))  severity failure;
	assert RAM(16745) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(16745))))  severity failure;
	assert RAM(16746) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(16746))))  severity failure;
	assert RAM(16747) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(16747))))  severity failure;
	assert RAM(16748) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(16748))))  severity failure;
	assert RAM(16749) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(16749))))  severity failure;
	assert RAM(16750) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(16750))))  severity failure;
	assert RAM(16751) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(16751))))  severity failure;
	assert RAM(16752) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(16752))))  severity failure;
	assert RAM(16753) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(16753))))  severity failure;
	assert RAM(16754) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(16754))))  severity failure;
	assert RAM(16755) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(16755))))  severity failure;
	assert RAM(16756) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(16756))))  severity failure;
	assert RAM(16757) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(16757))))  severity failure;
	assert RAM(16758) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(16758))))  severity failure;
	assert RAM(16759) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(16759))))  severity failure;
	assert RAM(16760) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(16760))))  severity failure;
	assert RAM(16761) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(16761))))  severity failure;
	assert RAM(16762) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(16762))))  severity failure;
	assert RAM(16763) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(16763))))  severity failure;
	assert RAM(16764) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(16764))))  severity failure;
	assert RAM(16765) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(16765))))  severity failure;
	assert RAM(16766) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(16766))))  severity failure;
	assert RAM(16767) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(16767))))  severity failure;
	assert RAM(16768) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(16768))))  severity failure;
	assert RAM(16769) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(16769))))  severity failure;
	assert RAM(16770) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(16770))))  severity failure;
	assert RAM(16771) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(16771))))  severity failure;
	assert RAM(16772) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(16772))))  severity failure;
	assert RAM(16773) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(16773))))  severity failure;
	assert RAM(16774) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(16774))))  severity failure;
	assert RAM(16775) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16775))))  severity failure;
	assert RAM(16776) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(16776))))  severity failure;
	assert RAM(16777) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(16777))))  severity failure;
	assert RAM(16778) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(16778))))  severity failure;
	assert RAM(16779) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(16779))))  severity failure;
	assert RAM(16780) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(16780))))  severity failure;
	assert RAM(16781) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(16781))))  severity failure;
	assert RAM(16782) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(16782))))  severity failure;
	assert RAM(16783) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16783))))  severity failure;
	assert RAM(16784) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(16784))))  severity failure;
	assert RAM(16785) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(16785))))  severity failure;
	assert RAM(16786) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(16786))))  severity failure;
	assert RAM(16787) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(16787))))  severity failure;
	assert RAM(16788) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(16788))))  severity failure;
	assert RAM(16789) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(16789))))  severity failure;
	assert RAM(16790) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(16790))))  severity failure;
	assert RAM(16791) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(16791))))  severity failure;
	assert RAM(16792) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(16792))))  severity failure;
	assert RAM(16793) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(16793))))  severity failure;
	assert RAM(16794) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(16794))))  severity failure;
	assert RAM(16795) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(16795))))  severity failure;
	assert RAM(16796) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(16796))))  severity failure;
	assert RAM(16797) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(16797))))  severity failure;
	assert RAM(16798) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(16798))))  severity failure;
	assert RAM(16799) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(16799))))  severity failure;
	assert RAM(16800) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(16800))))  severity failure;
	assert RAM(16801) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(16801))))  severity failure;
	assert RAM(16802) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(16802))))  severity failure;
	assert RAM(16803) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(16803))))  severity failure;
	assert RAM(16804) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(16804))))  severity failure;
	assert RAM(16805) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(16805))))  severity failure;
	assert RAM(16806) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(16806))))  severity failure;
	assert RAM(16807) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(16807))))  severity failure;
	assert RAM(16808) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16808))))  severity failure;
	assert RAM(16809) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(16809))))  severity failure;
	assert RAM(16810) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(16810))))  severity failure;
	assert RAM(16811) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(16811))))  severity failure;
	assert RAM(16812) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16812))))  severity failure;
	assert RAM(16813) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(16813))))  severity failure;
	assert RAM(16814) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(16814))))  severity failure;
	assert RAM(16815) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(16815))))  severity failure;
	assert RAM(16816) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(16816))))  severity failure;
	assert RAM(16817) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(16817))))  severity failure;
	assert RAM(16818) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(16818))))  severity failure;
	assert RAM(16819) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(16819))))  severity failure;
	assert RAM(16820) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16820))))  severity failure;
	assert RAM(16821) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(16821))))  severity failure;
	assert RAM(16822) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16822))))  severity failure;
	assert RAM(16823) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(16823))))  severity failure;
	assert RAM(16824) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(16824))))  severity failure;
	assert RAM(16825) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(16825))))  severity failure;
	assert RAM(16826) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16826))))  severity failure;
	assert RAM(16827) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(16827))))  severity failure;
	assert RAM(16828) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(16828))))  severity failure;
	assert RAM(16829) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(16829))))  severity failure;
	assert RAM(16830) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(16830))))  severity failure;
	assert RAM(16831) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(16831))))  severity failure;
	assert RAM(16832) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(16832))))  severity failure;
	assert RAM(16833) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(16833))))  severity failure;
	assert RAM(16834) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(16834))))  severity failure;
	assert RAM(16835) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(16835))))  severity failure;
	assert RAM(16836) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(16836))))  severity failure;
	assert RAM(16837) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(16837))))  severity failure;
	assert RAM(16838) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16838))))  severity failure;
	assert RAM(16839) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(16839))))  severity failure;
	assert RAM(16840) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16840))))  severity failure;
	assert RAM(16841) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(16841))))  severity failure;
	assert RAM(16842) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(16842))))  severity failure;
	assert RAM(16843) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16843))))  severity failure;
	assert RAM(16844) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16844))))  severity failure;
	assert RAM(16845) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(16845))))  severity failure;
	assert RAM(16846) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(16846))))  severity failure;
	assert RAM(16847) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16847))))  severity failure;
	assert RAM(16848) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(16848))))  severity failure;
	assert RAM(16849) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(16849))))  severity failure;
	assert RAM(16850) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(16850))))  severity failure;
	assert RAM(16851) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(16851))))  severity failure;
	assert RAM(16852) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(16852))))  severity failure;
	assert RAM(16853) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(16853))))  severity failure;
	assert RAM(16854) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(16854))))  severity failure;
	assert RAM(16855) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(16855))))  severity failure;
	assert RAM(16856) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(16856))))  severity failure;
	assert RAM(16857) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(16857))))  severity failure;
	assert RAM(16858) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(16858))))  severity failure;
	assert RAM(16859) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(16859))))  severity failure;
	assert RAM(16860) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(16860))))  severity failure;
	assert RAM(16861) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(16861))))  severity failure;
	assert RAM(16862) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(16862))))  severity failure;
	assert RAM(16863) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(16863))))  severity failure;
	assert RAM(16864) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(16864))))  severity failure;
	assert RAM(16865) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16865))))  severity failure;
	assert RAM(16866) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(16866))))  severity failure;
	assert RAM(16867) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(16867))))  severity failure;
	assert RAM(16868) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(16868))))  severity failure;
	assert RAM(16869) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16869))))  severity failure;
	assert RAM(16870) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(16870))))  severity failure;
	assert RAM(16871) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(16871))))  severity failure;
	assert RAM(16872) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(16872))))  severity failure;
	assert RAM(16873) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(16873))))  severity failure;
	assert RAM(16874) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(16874))))  severity failure;
	assert RAM(16875) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(16875))))  severity failure;
	assert RAM(16876) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(16876))))  severity failure;
	assert RAM(16877) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(16877))))  severity failure;
	assert RAM(16878) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(16878))))  severity failure;
	assert RAM(16879) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(16879))))  severity failure;
	assert RAM(16880) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(16880))))  severity failure;
	assert RAM(16881) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16881))))  severity failure;
	assert RAM(16882) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(16882))))  severity failure;
	assert RAM(16883) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(16883))))  severity failure;
	assert RAM(16884) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(16884))))  severity failure;
	assert RAM(16885) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(16885))))  severity failure;
	assert RAM(16886) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(16886))))  severity failure;
	assert RAM(16887) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(16887))))  severity failure;
	assert RAM(16888) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(16888))))  severity failure;
	assert RAM(16889) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(16889))))  severity failure;
	assert RAM(16890) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(16890))))  severity failure;
	assert RAM(16891) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(16891))))  severity failure;
	assert RAM(16892) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(16892))))  severity failure;
	assert RAM(16893) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(16893))))  severity failure;
	assert RAM(16894) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(16894))))  severity failure;
	assert RAM(16895) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16895))))  severity failure;
	assert RAM(16896) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16896))))  severity failure;
	assert RAM(16897) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(16897))))  severity failure;
	assert RAM(16898) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(16898))))  severity failure;
	assert RAM(16899) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(16899))))  severity failure;
	assert RAM(16900) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(16900))))  severity failure;
	assert RAM(16901) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(16901))))  severity failure;
	assert RAM(16902) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(16902))))  severity failure;
	assert RAM(16903) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(16903))))  severity failure;
	assert RAM(16904) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(16904))))  severity failure;
	assert RAM(16905) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(16905))))  severity failure;
	assert RAM(16906) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(16906))))  severity failure;
	assert RAM(16907) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(16907))))  severity failure;
	assert RAM(16908) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(16908))))  severity failure;
	assert RAM(16909) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(16909))))  severity failure;
	assert RAM(16910) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(16910))))  severity failure;
	assert RAM(16911) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(16911))))  severity failure;
	assert RAM(16912) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(16912))))  severity failure;
	assert RAM(16913) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(16913))))  severity failure;
	assert RAM(16914) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(16914))))  severity failure;
	assert RAM(16915) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(16915))))  severity failure;
	assert RAM(16916) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(16916))))  severity failure;
	assert RAM(16917) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(16917))))  severity failure;
	assert RAM(16918) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(16918))))  severity failure;
	assert RAM(16919) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(16919))))  severity failure;
	assert RAM(16920) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(16920))))  severity failure;
	assert RAM(16921) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(16921))))  severity failure;
	assert RAM(16922) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(16922))))  severity failure;
	assert RAM(16923) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(16923))))  severity failure;
	assert RAM(16924) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(16924))))  severity failure;
	assert RAM(16925) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(16925))))  severity failure;
	assert RAM(16926) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(16926))))  severity failure;
	assert RAM(16927) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(16927))))  severity failure;
	assert RAM(16928) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(16928))))  severity failure;
	assert RAM(16929) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(16929))))  severity failure;
	assert RAM(16930) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(16930))))  severity failure;
	assert RAM(16931) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(16931))))  severity failure;
	assert RAM(16932) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(16932))))  severity failure;
	assert RAM(16933) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(16933))))  severity failure;
	assert RAM(16934) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(16934))))  severity failure;
	assert RAM(16935) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(16935))))  severity failure;
	assert RAM(16936) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(16936))))  severity failure;
	assert RAM(16937) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16937))))  severity failure;
	assert RAM(16938) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(16938))))  severity failure;
	assert RAM(16939) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(16939))))  severity failure;
	assert RAM(16940) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(16940))))  severity failure;
	assert RAM(16941) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(16941))))  severity failure;
	assert RAM(16942) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(16942))))  severity failure;
	assert RAM(16943) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(16943))))  severity failure;
	assert RAM(16944) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(16944))))  severity failure;
	assert RAM(16945) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(16945))))  severity failure;
	assert RAM(16946) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(16946))))  severity failure;
	assert RAM(16947) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(16947))))  severity failure;
	assert RAM(16948) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(16948))))  severity failure;
	assert RAM(16949) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(16949))))  severity failure;
	assert RAM(16950) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(16950))))  severity failure;
	assert RAM(16951) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(16951))))  severity failure;
	assert RAM(16952) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(16952))))  severity failure;
	assert RAM(16953) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16953))))  severity failure;
	assert RAM(16954) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(16954))))  severity failure;
	assert RAM(16955) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(16955))))  severity failure;
	assert RAM(16956) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(16956))))  severity failure;
	assert RAM(16957) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(16957))))  severity failure;
	assert RAM(16958) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(16958))))  severity failure;
	assert RAM(16959) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(16959))))  severity failure;
	assert RAM(16960) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(16960))))  severity failure;
	assert RAM(16961) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(16961))))  severity failure;
	assert RAM(16962) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(16962))))  severity failure;
	assert RAM(16963) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(16963))))  severity failure;
	assert RAM(16964) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(16964))))  severity failure;
	assert RAM(16965) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(16965))))  severity failure;
	assert RAM(16966) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(16966))))  severity failure;
	assert RAM(16967) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(16967))))  severity failure;
	assert RAM(16968) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(16968))))  severity failure;
	assert RAM(16969) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(16969))))  severity failure;
	assert RAM(16970) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(16970))))  severity failure;
	assert RAM(16971) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(16971))))  severity failure;
	assert RAM(16972) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(16972))))  severity failure;
	assert RAM(16973) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(16973))))  severity failure;
	assert RAM(16974) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(16974))))  severity failure;
	assert RAM(16975) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(16975))))  severity failure;
	assert RAM(16976) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(16976))))  severity failure;
	assert RAM(16977) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(16977))))  severity failure;
	assert RAM(16978) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(16978))))  severity failure;
	assert RAM(16979) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(16979))))  severity failure;
	assert RAM(16980) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(16980))))  severity failure;
	assert RAM(16981) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(16981))))  severity failure;
	assert RAM(16982) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(16982))))  severity failure;
	assert RAM(16983) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(16983))))  severity failure;
	assert RAM(16984) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(16984))))  severity failure;
	assert RAM(16985) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(16985))))  severity failure;
	assert RAM(16986) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(16986))))  severity failure;
	assert RAM(16987) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(16987))))  severity failure;
	assert RAM(16988) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(16988))))  severity failure;
	assert RAM(16989) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(16989))))  severity failure;
	assert RAM(16990) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(16990))))  severity failure;
	assert RAM(16991) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(16991))))  severity failure;
	assert RAM(16992) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(16992))))  severity failure;
	assert RAM(16993) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(16993))))  severity failure;
	assert RAM(16994) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(16994))))  severity failure;
	assert RAM(16995) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(16995))))  severity failure;
	assert RAM(16996) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(16996))))  severity failure;
	assert RAM(16997) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(16997))))  severity failure;
	assert RAM(16998) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(16998))))  severity failure;
	assert RAM(16999) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(16999))))  severity failure;
	assert RAM(17000) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(17000))))  severity failure;
	assert RAM(17001) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(17001))))  severity failure;
	assert RAM(17002) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(17002))))  severity failure;
	assert RAM(17003) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(17003))))  severity failure;
	assert RAM(17004) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(17004))))  severity failure;
	assert RAM(17005) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17005))))  severity failure;
	assert RAM(17006) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(17006))))  severity failure;
	assert RAM(17007) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(17007))))  severity failure;
	assert RAM(17008) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(17008))))  severity failure;
	assert RAM(17009) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(17009))))  severity failure;
	assert RAM(17010) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(17010))))  severity failure;
	assert RAM(17011) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(17011))))  severity failure;
	assert RAM(17012) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(17012))))  severity failure;
	assert RAM(17013) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17013))))  severity failure;
	assert RAM(17014) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17014))))  severity failure;
	assert RAM(17015) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(17015))))  severity failure;
	assert RAM(17016) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(17016))))  severity failure;
	assert RAM(17017) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(17017))))  severity failure;
	assert RAM(17018) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17018))))  severity failure;
	assert RAM(17019) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17019))))  severity failure;
	assert RAM(17020) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17020))))  severity failure;
	assert RAM(17021) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17021))))  severity failure;
	assert RAM(17022) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(17022))))  severity failure;
	assert RAM(17023) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(17023))))  severity failure;
	assert RAM(17024) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(17024))))  severity failure;
	assert RAM(17025) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(17025))))  severity failure;
	assert RAM(17026) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(17026))))  severity failure;
	assert RAM(17027) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(17027))))  severity failure;
	assert RAM(17028) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17028))))  severity failure;
	assert RAM(17029) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(17029))))  severity failure;
	assert RAM(17030) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(17030))))  severity failure;
	assert RAM(17031) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17031))))  severity failure;
	assert RAM(17032) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(17032))))  severity failure;
	assert RAM(17033) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(17033))))  severity failure;
	assert RAM(17034) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17034))))  severity failure;
	assert RAM(17035) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17035))))  severity failure;
	assert RAM(17036) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(17036))))  severity failure;
	assert RAM(17037) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(17037))))  severity failure;
	assert RAM(17038) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(17038))))  severity failure;
	assert RAM(17039) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(17039))))  severity failure;
	assert RAM(17040) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(17040))))  severity failure;
	assert RAM(17041) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17041))))  severity failure;
	assert RAM(17042) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(17042))))  severity failure;
	assert RAM(17043) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(17043))))  severity failure;
	assert RAM(17044) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(17044))))  severity failure;
	assert RAM(17045) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(17045))))  severity failure;
	assert RAM(17046) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(17046))))  severity failure;
	assert RAM(17047) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17047))))  severity failure;
	assert RAM(17048) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(17048))))  severity failure;
	assert RAM(17049) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17049))))  severity failure;
	assert RAM(17050) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(17050))))  severity failure;
	assert RAM(17051) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(17051))))  severity failure;
	assert RAM(17052) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17052))))  severity failure;
	assert RAM(17053) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17053))))  severity failure;
	assert RAM(17054) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17054))))  severity failure;
	assert RAM(17055) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(17055))))  severity failure;
	assert RAM(17056) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(17056))))  severity failure;
	assert RAM(17057) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(17057))))  severity failure;
	assert RAM(17058) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(17058))))  severity failure;
	assert RAM(17059) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(17059))))  severity failure;
	assert RAM(17060) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(17060))))  severity failure;
	assert RAM(17061) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(17061))))  severity failure;
	assert RAM(17062) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(17062))))  severity failure;
	assert RAM(17063) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(17063))))  severity failure;
	assert RAM(17064) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(17064))))  severity failure;
	assert RAM(17065) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(17065))))  severity failure;
	assert RAM(17066) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(17066))))  severity failure;
	assert RAM(17067) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(17067))))  severity failure;
	assert RAM(17068) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(17068))))  severity failure;
	assert RAM(17069) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(17069))))  severity failure;
	assert RAM(17070) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(17070))))  severity failure;
	assert RAM(17071) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17071))))  severity failure;
	assert RAM(17072) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(17072))))  severity failure;
	assert RAM(17073) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(17073))))  severity failure;
	assert RAM(17074) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17074))))  severity failure;
	assert RAM(17075) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(17075))))  severity failure;
	assert RAM(17076) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(17076))))  severity failure;
	assert RAM(17077) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17077))))  severity failure;
	assert RAM(17078) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(17078))))  severity failure;
	assert RAM(17079) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(17079))))  severity failure;
	assert RAM(17080) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(17080))))  severity failure;
	assert RAM(17081) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17081))))  severity failure;
	assert RAM(17082) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17082))))  severity failure;
	assert RAM(17083) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(17083))))  severity failure;
	assert RAM(17084) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(17084))))  severity failure;
	assert RAM(17085) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17085))))  severity failure;
	assert RAM(17086) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17086))))  severity failure;
	assert RAM(17087) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(17087))))  severity failure;
	assert RAM(17088) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(17088))))  severity failure;
	assert RAM(17089) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17089))))  severity failure;
	assert RAM(17090) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17090))))  severity failure;
	assert RAM(17091) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(17091))))  severity failure;
	assert RAM(17092) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(17092))))  severity failure;
	assert RAM(17093) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17093))))  severity failure;
	assert RAM(17094) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(17094))))  severity failure;
	assert RAM(17095) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(17095))))  severity failure;
	assert RAM(17096) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(17096))))  severity failure;
	assert RAM(17097) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(17097))))  severity failure;
	assert RAM(17098) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(17098))))  severity failure;
	assert RAM(17099) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(17099))))  severity failure;
	assert RAM(17100) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(17100))))  severity failure;
	assert RAM(17101) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(17101))))  severity failure;
	assert RAM(17102) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17102))))  severity failure;
	assert RAM(17103) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17103))))  severity failure;
	assert RAM(17104) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17104))))  severity failure;
	assert RAM(17105) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17105))))  severity failure;
	assert RAM(17106) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17106))))  severity failure;
	assert RAM(17107) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(17107))))  severity failure;
	assert RAM(17108) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(17108))))  severity failure;
	assert RAM(17109) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(17109))))  severity failure;
	assert RAM(17110) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(17110))))  severity failure;
	assert RAM(17111) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(17111))))  severity failure;
	assert RAM(17112) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(17112))))  severity failure;
	assert RAM(17113) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(17113))))  severity failure;
	assert RAM(17114) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(17114))))  severity failure;
	assert RAM(17115) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(17115))))  severity failure;
	assert RAM(17116) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(17116))))  severity failure;
	assert RAM(17117) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(17117))))  severity failure;
	assert RAM(17118) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17118))))  severity failure;
	assert RAM(17119) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(17119))))  severity failure;
	assert RAM(17120) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(17120))))  severity failure;
	assert RAM(17121) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(17121))))  severity failure;
	assert RAM(17122) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(17122))))  severity failure;
	assert RAM(17123) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(17123))))  severity failure;
	assert RAM(17124) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17124))))  severity failure;
	assert RAM(17125) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(17125))))  severity failure;
	assert RAM(17126) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(17126))))  severity failure;
	assert RAM(17127) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(17127))))  severity failure;
	assert RAM(17128) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(17128))))  severity failure;
	assert RAM(17129) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(17129))))  severity failure;
	assert RAM(17130) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(17130))))  severity failure;
	assert RAM(17131) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17131))))  severity failure;
	assert RAM(17132) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(17132))))  severity failure;
	assert RAM(17133) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(17133))))  severity failure;
	assert RAM(17134) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(17134))))  severity failure;
	assert RAM(17135) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17135))))  severity failure;
	assert RAM(17136) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(17136))))  severity failure;
	assert RAM(17137) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(17137))))  severity failure;
	assert RAM(17138) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17138))))  severity failure;
	assert RAM(17139) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(17139))))  severity failure;
	assert RAM(17140) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(17140))))  severity failure;
	assert RAM(17141) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(17141))))  severity failure;
	assert RAM(17142) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(17142))))  severity failure;
	assert RAM(17143) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17143))))  severity failure;
	assert RAM(17144) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(17144))))  severity failure;
	assert RAM(17145) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17145))))  severity failure;
	assert RAM(17146) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(17146))))  severity failure;
	assert RAM(17147) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(17147))))  severity failure;
	assert RAM(17148) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17148))))  severity failure;
	assert RAM(17149) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(17149))))  severity failure;
	assert RAM(17150) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(17150))))  severity failure;
	assert RAM(17151) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(17151))))  severity failure;
	assert RAM(17152) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17152))))  severity failure;
	assert RAM(17153) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17153))))  severity failure;
	assert RAM(17154) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(17154))))  severity failure;
	assert RAM(17155) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17155))))  severity failure;
	assert RAM(17156) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(17156))))  severity failure;
	assert RAM(17157) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(17157))))  severity failure;
	assert RAM(17158) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17158))))  severity failure;
	assert RAM(17159) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(17159))))  severity failure;
	assert RAM(17160) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17160))))  severity failure;
	assert RAM(17161) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(17161))))  severity failure;
	assert RAM(17162) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17162))))  severity failure;
	assert RAM(17163) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17163))))  severity failure;
	assert RAM(17164) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(17164))))  severity failure;
	assert RAM(17165) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(17165))))  severity failure;
	assert RAM(17166) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(17166))))  severity failure;
	assert RAM(17167) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(17167))))  severity failure;
	assert RAM(17168) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(17168))))  severity failure;
	assert RAM(17169) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(17169))))  severity failure;
	assert RAM(17170) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(17170))))  severity failure;
	assert RAM(17171) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(17171))))  severity failure;
	assert RAM(17172) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(17172))))  severity failure;
	assert RAM(17173) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17173))))  severity failure;
	assert RAM(17174) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(17174))))  severity failure;
	assert RAM(17175) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(17175))))  severity failure;
	assert RAM(17176) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(17176))))  severity failure;
	assert RAM(17177) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17177))))  severity failure;
	assert RAM(17178) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17178))))  severity failure;
	assert RAM(17179) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17179))))  severity failure;
	assert RAM(17180) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(17180))))  severity failure;
	assert RAM(17181) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(17181))))  severity failure;
	assert RAM(17182) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(17182))))  severity failure;
	assert RAM(17183) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(17183))))  severity failure;
	assert RAM(17184) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(17184))))  severity failure;
	assert RAM(17185) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(17185))))  severity failure;
	assert RAM(17186) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(17186))))  severity failure;
	assert RAM(17187) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(17187))))  severity failure;
	assert RAM(17188) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(17188))))  severity failure;
	assert RAM(17189) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(17189))))  severity failure;
	assert RAM(17190) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(17190))))  severity failure;
	assert RAM(17191) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(17191))))  severity failure;
	assert RAM(17192) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(17192))))  severity failure;
	assert RAM(17193) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(17193))))  severity failure;
	assert RAM(17194) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(17194))))  severity failure;
	assert RAM(17195) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(17195))))  severity failure;
	assert RAM(17196) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(17196))))  severity failure;
	assert RAM(17197) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(17197))))  severity failure;
	assert RAM(17198) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(17198))))  severity failure;
	assert RAM(17199) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17199))))  severity failure;
	assert RAM(17200) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(17200))))  severity failure;
	assert RAM(17201) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(17201))))  severity failure;
	assert RAM(17202) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(17202))))  severity failure;
	assert RAM(17203) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(17203))))  severity failure;
	assert RAM(17204) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(17204))))  severity failure;
	assert RAM(17205) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17205))))  severity failure;
	assert RAM(17206) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(17206))))  severity failure;
	assert RAM(17207) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(17207))))  severity failure;
	assert RAM(17208) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17208))))  severity failure;
	assert RAM(17209) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(17209))))  severity failure;
	assert RAM(17210) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(17210))))  severity failure;
	assert RAM(17211) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(17211))))  severity failure;
	assert RAM(17212) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17212))))  severity failure;
	assert RAM(17213) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17213))))  severity failure;
	assert RAM(17214) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(17214))))  severity failure;
	assert RAM(17215) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(17215))))  severity failure;
	assert RAM(17216) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(17216))))  severity failure;
	assert RAM(17217) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(17217))))  severity failure;
	assert RAM(17218) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(17218))))  severity failure;
	assert RAM(17219) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17219))))  severity failure;
	assert RAM(17220) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(17220))))  severity failure;
	assert RAM(17221) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(17221))))  severity failure;
	assert RAM(17222) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(17222))))  severity failure;
	assert RAM(17223) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17223))))  severity failure;
	assert RAM(17224) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(17224))))  severity failure;
	assert RAM(17225) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(17225))))  severity failure;
	assert RAM(17226) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(17226))))  severity failure;
	assert RAM(17227) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17227))))  severity failure;
	assert RAM(17228) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(17228))))  severity failure;
	assert RAM(17229) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17229))))  severity failure;
	assert RAM(17230) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17230))))  severity failure;
	assert RAM(17231) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17231))))  severity failure;
	assert RAM(17232) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17232))))  severity failure;
	assert RAM(17233) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(17233))))  severity failure;
	assert RAM(17234) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(17234))))  severity failure;
	assert RAM(17235) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(17235))))  severity failure;
	assert RAM(17236) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(17236))))  severity failure;
	assert RAM(17237) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(17237))))  severity failure;
	assert RAM(17238) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(17238))))  severity failure;
	assert RAM(17239) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(17239))))  severity failure;
	assert RAM(17240) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(17240))))  severity failure;
	assert RAM(17241) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(17241))))  severity failure;
	assert RAM(17242) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17242))))  severity failure;
	assert RAM(17243) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(17243))))  severity failure;
	assert RAM(17244) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(17244))))  severity failure;
	assert RAM(17245) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(17245))))  severity failure;
	assert RAM(17246) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17246))))  severity failure;
	assert RAM(17247) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(17247))))  severity failure;
	assert RAM(17248) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(17248))))  severity failure;
	assert RAM(17249) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(17249))))  severity failure;
	assert RAM(17250) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(17250))))  severity failure;
	assert RAM(17251) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17251))))  severity failure;
	assert RAM(17252) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(17252))))  severity failure;
	assert RAM(17253) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(17253))))  severity failure;
	assert RAM(17254) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(17254))))  severity failure;
	assert RAM(17255) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(17255))))  severity failure;
	assert RAM(17256) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17256))))  severity failure;
	assert RAM(17257) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(17257))))  severity failure;
	assert RAM(17258) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(17258))))  severity failure;
	assert RAM(17259) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17259))))  severity failure;
	assert RAM(17260) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17260))))  severity failure;
	assert RAM(17261) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17261))))  severity failure;
	assert RAM(17262) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(17262))))  severity failure;
	assert RAM(17263) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17263))))  severity failure;
	assert RAM(17264) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17264))))  severity failure;
	assert RAM(17265) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(17265))))  severity failure;
	assert RAM(17266) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(17266))))  severity failure;
	assert RAM(17267) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(17267))))  severity failure;
	assert RAM(17268) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(17268))))  severity failure;
	assert RAM(17269) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(17269))))  severity failure;
	assert RAM(17270) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17270))))  severity failure;
	assert RAM(17271) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17271))))  severity failure;
	assert RAM(17272) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17272))))  severity failure;
	assert RAM(17273) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(17273))))  severity failure;
	assert RAM(17274) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17274))))  severity failure;
	assert RAM(17275) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17275))))  severity failure;
	assert RAM(17276) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(17276))))  severity failure;
	assert RAM(17277) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(17277))))  severity failure;
	assert RAM(17278) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(17278))))  severity failure;
	assert RAM(17279) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(17279))))  severity failure;
	assert RAM(17280) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17280))))  severity failure;
	assert RAM(17281) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(17281))))  severity failure;
	assert RAM(17282) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(17282))))  severity failure;
	assert RAM(17283) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(17283))))  severity failure;
	assert RAM(17284) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17284))))  severity failure;
	assert RAM(17285) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(17285))))  severity failure;
	assert RAM(17286) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17286))))  severity failure;
	assert RAM(17287) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(17287))))  severity failure;
	assert RAM(17288) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(17288))))  severity failure;
	assert RAM(17289) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(17289))))  severity failure;
	assert RAM(17290) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17290))))  severity failure;
	assert RAM(17291) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(17291))))  severity failure;
	assert RAM(17292) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(17292))))  severity failure;
	assert RAM(17293) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(17293))))  severity failure;
	assert RAM(17294) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17294))))  severity failure;
	assert RAM(17295) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(17295))))  severity failure;
	assert RAM(17296) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17296))))  severity failure;
	assert RAM(17297) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(17297))))  severity failure;
	assert RAM(17298) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(17298))))  severity failure;
	assert RAM(17299) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(17299))))  severity failure;
	assert RAM(17300) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(17300))))  severity failure;
	assert RAM(17301) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17301))))  severity failure;
	assert RAM(17302) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(17302))))  severity failure;
	assert RAM(17303) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(17303))))  severity failure;
	assert RAM(17304) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17304))))  severity failure;
	assert RAM(17305) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(17305))))  severity failure;
	assert RAM(17306) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(17306))))  severity failure;
	assert RAM(17307) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17307))))  severity failure;
	assert RAM(17308) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(17308))))  severity failure;
	assert RAM(17309) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(17309))))  severity failure;
	assert RAM(17310) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(17310))))  severity failure;
	assert RAM(17311) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(17311))))  severity failure;
	assert RAM(17312) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(17312))))  severity failure;
	assert RAM(17313) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(17313))))  severity failure;
	assert RAM(17314) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(17314))))  severity failure;
	assert RAM(17315) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(17315))))  severity failure;
	assert RAM(17316) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17316))))  severity failure;
	assert RAM(17317) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17317))))  severity failure;
	assert RAM(17318) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(17318))))  severity failure;
	assert RAM(17319) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(17319))))  severity failure;
	assert RAM(17320) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(17320))))  severity failure;
	assert RAM(17321) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17321))))  severity failure;
	assert RAM(17322) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(17322))))  severity failure;
	assert RAM(17323) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(17323))))  severity failure;
	assert RAM(17324) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17324))))  severity failure;
	assert RAM(17325) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(17325))))  severity failure;
	assert RAM(17326) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(17326))))  severity failure;
	assert RAM(17327) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(17327))))  severity failure;
	assert RAM(17328) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17328))))  severity failure;
	assert RAM(17329) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(17329))))  severity failure;
	assert RAM(17330) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(17330))))  severity failure;
	assert RAM(17331) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(17331))))  severity failure;
	assert RAM(17332) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(17332))))  severity failure;
	assert RAM(17333) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17333))))  severity failure;
	assert RAM(17334) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(17334))))  severity failure;
	assert RAM(17335) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(17335))))  severity failure;
	assert RAM(17336) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(17336))))  severity failure;
	assert RAM(17337) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(17337))))  severity failure;
	assert RAM(17338) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(17338))))  severity failure;
	assert RAM(17339) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(17339))))  severity failure;
	assert RAM(17340) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17340))))  severity failure;
	assert RAM(17341) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17341))))  severity failure;
	assert RAM(17342) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(17342))))  severity failure;
	assert RAM(17343) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(17343))))  severity failure;
	assert RAM(17344) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(17344))))  severity failure;
	assert RAM(17345) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17345))))  severity failure;
	assert RAM(17346) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(17346))))  severity failure;
	assert RAM(17347) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(17347))))  severity failure;
	assert RAM(17348) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(17348))))  severity failure;
	assert RAM(17349) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(17349))))  severity failure;
	assert RAM(17350) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(17350))))  severity failure;
	assert RAM(17351) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(17351))))  severity failure;
	assert RAM(17352) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(17352))))  severity failure;
	assert RAM(17353) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(17353))))  severity failure;
	assert RAM(17354) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(17354))))  severity failure;
	assert RAM(17355) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(17355))))  severity failure;
	assert RAM(17356) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(17356))))  severity failure;
	assert RAM(17357) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17357))))  severity failure;
	assert RAM(17358) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17358))))  severity failure;
	assert RAM(17359) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17359))))  severity failure;
	assert RAM(17360) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17360))))  severity failure;
	assert RAM(17361) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(17361))))  severity failure;
	assert RAM(17362) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(17362))))  severity failure;
	assert RAM(17363) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17363))))  severity failure;
	assert RAM(17364) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(17364))))  severity failure;
	assert RAM(17365) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(17365))))  severity failure;
	assert RAM(17366) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(17366))))  severity failure;
	assert RAM(17367) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(17367))))  severity failure;
	assert RAM(17368) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17368))))  severity failure;
	assert RAM(17369) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(17369))))  severity failure;
	assert RAM(17370) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(17370))))  severity failure;
	assert RAM(17371) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(17371))))  severity failure;
	assert RAM(17372) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(17372))))  severity failure;
	assert RAM(17373) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(17373))))  severity failure;
	assert RAM(17374) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(17374))))  severity failure;
	assert RAM(17375) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(17375))))  severity failure;
	assert RAM(17376) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17376))))  severity failure;
	assert RAM(17377) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(17377))))  severity failure;
	assert RAM(17378) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(17378))))  severity failure;
	assert RAM(17379) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(17379))))  severity failure;
	assert RAM(17380) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(17380))))  severity failure;
	assert RAM(17381) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(17381))))  severity failure;
	assert RAM(17382) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(17382))))  severity failure;
	assert RAM(17383) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(17383))))  severity failure;
	assert RAM(17384) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(17384))))  severity failure;
	assert RAM(17385) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(17385))))  severity failure;
	assert RAM(17386) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(17386))))  severity failure;
	assert RAM(17387) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(17387))))  severity failure;
	assert RAM(17388) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(17388))))  severity failure;
	assert RAM(17389) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(17389))))  severity failure;
	assert RAM(17390) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17390))))  severity failure;
	assert RAM(17391) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(17391))))  severity failure;
	assert RAM(17392) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(17392))))  severity failure;
	assert RAM(17393) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(17393))))  severity failure;
	assert RAM(17394) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(17394))))  severity failure;
	assert RAM(17395) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(17395))))  severity failure;
	assert RAM(17396) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(17396))))  severity failure;
	assert RAM(17397) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(17397))))  severity failure;
	assert RAM(17398) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(17398))))  severity failure;
	assert RAM(17399) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17399))))  severity failure;
	assert RAM(17400) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(17400))))  severity failure;
	assert RAM(17401) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17401))))  severity failure;
	assert RAM(17402) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(17402))))  severity failure;
	assert RAM(17403) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(17403))))  severity failure;
	assert RAM(17404) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(17404))))  severity failure;
	assert RAM(17405) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(17405))))  severity failure;
	assert RAM(17406) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17406))))  severity failure;
	assert RAM(17407) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(17407))))  severity failure;
	assert RAM(17408) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17408))))  severity failure;
	assert RAM(17409) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(17409))))  severity failure;
	assert RAM(17410) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(17410))))  severity failure;
	assert RAM(17411) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(17411))))  severity failure;
	assert RAM(17412) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(17412))))  severity failure;
	assert RAM(17413) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(17413))))  severity failure;
	assert RAM(17414) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(17414))))  severity failure;
	assert RAM(17415) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(17415))))  severity failure;
	assert RAM(17416) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(17416))))  severity failure;
	assert RAM(17417) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17417))))  severity failure;
	assert RAM(17418) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(17418))))  severity failure;
	assert RAM(17419) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(17419))))  severity failure;
	assert RAM(17420) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17420))))  severity failure;
	assert RAM(17421) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(17421))))  severity failure;
	assert RAM(17422) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(17422))))  severity failure;
	assert RAM(17423) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(17423))))  severity failure;
	assert RAM(17424) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17424))))  severity failure;
	assert RAM(17425) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(17425))))  severity failure;
	assert RAM(17426) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17426))))  severity failure;
	assert RAM(17427) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(17427))))  severity failure;
	assert RAM(17428) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(17428))))  severity failure;
	assert RAM(17429) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17429))))  severity failure;
	assert RAM(17430) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(17430))))  severity failure;
	assert RAM(17431) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17431))))  severity failure;
	assert RAM(17432) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17432))))  severity failure;
	assert RAM(17433) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17433))))  severity failure;
	assert RAM(17434) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17434))))  severity failure;
	assert RAM(17435) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17435))))  severity failure;
	assert RAM(17436) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17436))))  severity failure;
	assert RAM(17437) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(17437))))  severity failure;
	assert RAM(17438) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17438))))  severity failure;
	assert RAM(17439) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(17439))))  severity failure;
	assert RAM(17440) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(17440))))  severity failure;
	assert RAM(17441) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17441))))  severity failure;
	assert RAM(17442) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17442))))  severity failure;
	assert RAM(17443) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(17443))))  severity failure;
	assert RAM(17444) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17444))))  severity failure;
	assert RAM(17445) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17445))))  severity failure;
	assert RAM(17446) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(17446))))  severity failure;
	assert RAM(17447) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(17447))))  severity failure;
	assert RAM(17448) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17448))))  severity failure;
	assert RAM(17449) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(17449))))  severity failure;
	assert RAM(17450) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(17450))))  severity failure;
	assert RAM(17451) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(17451))))  severity failure;
	assert RAM(17452) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(17452))))  severity failure;
	assert RAM(17453) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17453))))  severity failure;
	assert RAM(17454) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(17454))))  severity failure;
	assert RAM(17455) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(17455))))  severity failure;
	assert RAM(17456) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(17456))))  severity failure;
	assert RAM(17457) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(17457))))  severity failure;
	assert RAM(17458) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(17458))))  severity failure;
	assert RAM(17459) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17459))))  severity failure;
	assert RAM(17460) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(17460))))  severity failure;
	assert RAM(17461) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(17461))))  severity failure;
	assert RAM(17462) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(17462))))  severity failure;
	assert RAM(17463) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(17463))))  severity failure;
	assert RAM(17464) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(17464))))  severity failure;
	assert RAM(17465) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(17465))))  severity failure;
	assert RAM(17466) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(17466))))  severity failure;
	assert RAM(17467) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(17467))))  severity failure;
	assert RAM(17468) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17468))))  severity failure;
	assert RAM(17469) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17469))))  severity failure;
	assert RAM(17470) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17470))))  severity failure;
	assert RAM(17471) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(17471))))  severity failure;
	assert RAM(17472) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(17472))))  severity failure;
	assert RAM(17473) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17473))))  severity failure;
	assert RAM(17474) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(17474))))  severity failure;
	assert RAM(17475) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(17475))))  severity failure;
	assert RAM(17476) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(17476))))  severity failure;
	assert RAM(17477) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(17477))))  severity failure;
	assert RAM(17478) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(17478))))  severity failure;
	assert RAM(17479) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(17479))))  severity failure;
	assert RAM(17480) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(17480))))  severity failure;
	assert RAM(17481) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(17481))))  severity failure;
	assert RAM(17482) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(17482))))  severity failure;
	assert RAM(17483) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17483))))  severity failure;
	assert RAM(17484) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(17484))))  severity failure;
	assert RAM(17485) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17485))))  severity failure;
	assert RAM(17486) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(17486))))  severity failure;
	assert RAM(17487) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(17487))))  severity failure;
	assert RAM(17488) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17488))))  severity failure;
	assert RAM(17489) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(17489))))  severity failure;
	assert RAM(17490) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17490))))  severity failure;
	assert RAM(17491) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17491))))  severity failure;
	assert RAM(17492) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(17492))))  severity failure;
	assert RAM(17493) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(17493))))  severity failure;
	assert RAM(17494) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17494))))  severity failure;
	assert RAM(17495) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(17495))))  severity failure;
	assert RAM(17496) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(17496))))  severity failure;
	assert RAM(17497) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(17497))))  severity failure;
	assert RAM(17498) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17498))))  severity failure;
	assert RAM(17499) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(17499))))  severity failure;
	assert RAM(17500) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17500))))  severity failure;
	assert RAM(17501) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(17501))))  severity failure;
	assert RAM(17502) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(17502))))  severity failure;
	assert RAM(17503) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(17503))))  severity failure;
	assert RAM(17504) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(17504))))  severity failure;
	assert RAM(17505) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(17505))))  severity failure;
	assert RAM(17506) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(17506))))  severity failure;
	assert RAM(17507) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17507))))  severity failure;
	assert RAM(17508) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(17508))))  severity failure;
	assert RAM(17509) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(17509))))  severity failure;
	assert RAM(17510) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(17510))))  severity failure;
	assert RAM(17511) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(17511))))  severity failure;
	assert RAM(17512) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(17512))))  severity failure;
	assert RAM(17513) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(17513))))  severity failure;
	assert RAM(17514) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(17514))))  severity failure;
	assert RAM(17515) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17515))))  severity failure;
	assert RAM(17516) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17516))))  severity failure;
	assert RAM(17517) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(17517))))  severity failure;
	assert RAM(17518) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17518))))  severity failure;
	assert RAM(17519) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(17519))))  severity failure;
	assert RAM(17520) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(17520))))  severity failure;
	assert RAM(17521) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17521))))  severity failure;
	assert RAM(17522) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(17522))))  severity failure;
	assert RAM(17523) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(17523))))  severity failure;
	assert RAM(17524) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17524))))  severity failure;
	assert RAM(17525) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17525))))  severity failure;
	assert RAM(17526) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(17526))))  severity failure;
	assert RAM(17527) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(17527))))  severity failure;
	assert RAM(17528) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17528))))  severity failure;
	assert RAM(17529) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(17529))))  severity failure;
	assert RAM(17530) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17530))))  severity failure;
	assert RAM(17531) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(17531))))  severity failure;
	assert RAM(17532) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17532))))  severity failure;
	assert RAM(17533) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(17533))))  severity failure;
	assert RAM(17534) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(17534))))  severity failure;
	assert RAM(17535) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17535))))  severity failure;
	assert RAM(17536) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(17536))))  severity failure;
	assert RAM(17537) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17537))))  severity failure;
	assert RAM(17538) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(17538))))  severity failure;
	assert RAM(17539) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17539))))  severity failure;
	assert RAM(17540) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(17540))))  severity failure;
	assert RAM(17541) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17541))))  severity failure;
	assert RAM(17542) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(17542))))  severity failure;
	assert RAM(17543) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17543))))  severity failure;
	assert RAM(17544) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17544))))  severity failure;
	assert RAM(17545) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(17545))))  severity failure;
	assert RAM(17546) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(17546))))  severity failure;
	assert RAM(17547) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(17547))))  severity failure;
	assert RAM(17548) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(17548))))  severity failure;
	assert RAM(17549) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17549))))  severity failure;
	assert RAM(17550) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17550))))  severity failure;
	assert RAM(17551) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17551))))  severity failure;
	assert RAM(17552) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17552))))  severity failure;
	assert RAM(17553) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(17553))))  severity failure;
	assert RAM(17554) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(17554))))  severity failure;
	assert RAM(17555) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(17555))))  severity failure;
	assert RAM(17556) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(17556))))  severity failure;
	assert RAM(17557) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(17557))))  severity failure;
	assert RAM(17558) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(17558))))  severity failure;
	assert RAM(17559) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17559))))  severity failure;
	assert RAM(17560) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17560))))  severity failure;
	assert RAM(17561) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(17561))))  severity failure;
	assert RAM(17562) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(17562))))  severity failure;
	assert RAM(17563) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17563))))  severity failure;
	assert RAM(17564) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(17564))))  severity failure;
	assert RAM(17565) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(17565))))  severity failure;
	assert RAM(17566) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(17566))))  severity failure;
	assert RAM(17567) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(17567))))  severity failure;
	assert RAM(17568) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(17568))))  severity failure;
	assert RAM(17569) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17569))))  severity failure;
	assert RAM(17570) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17570))))  severity failure;
	assert RAM(17571) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(17571))))  severity failure;
	assert RAM(17572) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(17572))))  severity failure;
	assert RAM(17573) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(17573))))  severity failure;
	assert RAM(17574) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(17574))))  severity failure;
	assert RAM(17575) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(17575))))  severity failure;
	assert RAM(17576) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17576))))  severity failure;
	assert RAM(17577) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(17577))))  severity failure;
	assert RAM(17578) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17578))))  severity failure;
	assert RAM(17579) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(17579))))  severity failure;
	assert RAM(17580) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17580))))  severity failure;
	assert RAM(17581) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(17581))))  severity failure;
	assert RAM(17582) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(17582))))  severity failure;
	assert RAM(17583) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(17583))))  severity failure;
	assert RAM(17584) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(17584))))  severity failure;
	assert RAM(17585) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(17585))))  severity failure;
	assert RAM(17586) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(17586))))  severity failure;
	assert RAM(17587) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17587))))  severity failure;
	assert RAM(17588) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(17588))))  severity failure;
	assert RAM(17589) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(17589))))  severity failure;
	assert RAM(17590) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(17590))))  severity failure;
	assert RAM(17591) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17591))))  severity failure;
	assert RAM(17592) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(17592))))  severity failure;
	assert RAM(17593) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17593))))  severity failure;
	assert RAM(17594) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(17594))))  severity failure;
	assert RAM(17595) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17595))))  severity failure;
	assert RAM(17596) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(17596))))  severity failure;
	assert RAM(17597) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17597))))  severity failure;
	assert RAM(17598) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(17598))))  severity failure;
	assert RAM(17599) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(17599))))  severity failure;
	assert RAM(17600) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(17600))))  severity failure;
	assert RAM(17601) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(17601))))  severity failure;
	assert RAM(17602) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(17602))))  severity failure;
	assert RAM(17603) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(17603))))  severity failure;
	assert RAM(17604) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(17604))))  severity failure;
	assert RAM(17605) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17605))))  severity failure;
	assert RAM(17606) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17606))))  severity failure;
	assert RAM(17607) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(17607))))  severity failure;
	assert RAM(17608) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(17608))))  severity failure;
	assert RAM(17609) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17609))))  severity failure;
	assert RAM(17610) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(17610))))  severity failure;
	assert RAM(17611) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(17611))))  severity failure;
	assert RAM(17612) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17612))))  severity failure;
	assert RAM(17613) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(17613))))  severity failure;
	assert RAM(17614) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17614))))  severity failure;
	assert RAM(17615) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(17615))))  severity failure;
	assert RAM(17616) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(17616))))  severity failure;
	assert RAM(17617) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(17617))))  severity failure;
	assert RAM(17618) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(17618))))  severity failure;
	assert RAM(17619) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17619))))  severity failure;
	assert RAM(17620) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(17620))))  severity failure;
	assert RAM(17621) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(17621))))  severity failure;
	assert RAM(17622) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(17622))))  severity failure;
	assert RAM(17623) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(17623))))  severity failure;
	assert RAM(17624) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(17624))))  severity failure;
	assert RAM(17625) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(17625))))  severity failure;
	assert RAM(17626) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(17626))))  severity failure;
	assert RAM(17627) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17627))))  severity failure;
	assert RAM(17628) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(17628))))  severity failure;
	assert RAM(17629) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(17629))))  severity failure;
	assert RAM(17630) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(17630))))  severity failure;
	assert RAM(17631) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(17631))))  severity failure;
	assert RAM(17632) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(17632))))  severity failure;
	assert RAM(17633) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(17633))))  severity failure;
	assert RAM(17634) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17634))))  severity failure;
	assert RAM(17635) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17635))))  severity failure;
	assert RAM(17636) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(17636))))  severity failure;
	assert RAM(17637) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(17637))))  severity failure;
	assert RAM(17638) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17638))))  severity failure;
	assert RAM(17639) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(17639))))  severity failure;
	assert RAM(17640) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(17640))))  severity failure;
	assert RAM(17641) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(17641))))  severity failure;
	assert RAM(17642) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17642))))  severity failure;
	assert RAM(17643) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17643))))  severity failure;
	assert RAM(17644) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17644))))  severity failure;
	assert RAM(17645) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(17645))))  severity failure;
	assert RAM(17646) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(17646))))  severity failure;
	assert RAM(17647) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(17647))))  severity failure;
	assert RAM(17648) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(17648))))  severity failure;
	assert RAM(17649) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(17649))))  severity failure;
	assert RAM(17650) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(17650))))  severity failure;
	assert RAM(17651) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(17651))))  severity failure;
	assert RAM(17652) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17652))))  severity failure;
	assert RAM(17653) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(17653))))  severity failure;
	assert RAM(17654) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(17654))))  severity failure;
	assert RAM(17655) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(17655))))  severity failure;
	assert RAM(17656) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17656))))  severity failure;
	assert RAM(17657) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(17657))))  severity failure;
	assert RAM(17658) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(17658))))  severity failure;
	assert RAM(17659) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17659))))  severity failure;
	assert RAM(17660) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17660))))  severity failure;
	assert RAM(17661) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(17661))))  severity failure;
	assert RAM(17662) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17662))))  severity failure;
	assert RAM(17663) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(17663))))  severity failure;
	assert RAM(17664) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(17664))))  severity failure;
	assert RAM(17665) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(17665))))  severity failure;
	assert RAM(17666) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(17666))))  severity failure;
	assert RAM(17667) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17667))))  severity failure;
	assert RAM(17668) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(17668))))  severity failure;
	assert RAM(17669) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(17669))))  severity failure;
	assert RAM(17670) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17670))))  severity failure;
	assert RAM(17671) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(17671))))  severity failure;
	assert RAM(17672) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(17672))))  severity failure;
	assert RAM(17673) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(17673))))  severity failure;
	assert RAM(17674) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17674))))  severity failure;
	assert RAM(17675) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(17675))))  severity failure;
	assert RAM(17676) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(17676))))  severity failure;
	assert RAM(17677) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(17677))))  severity failure;
	assert RAM(17678) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(17678))))  severity failure;
	assert RAM(17679) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(17679))))  severity failure;
	assert RAM(17680) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(17680))))  severity failure;
	assert RAM(17681) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(17681))))  severity failure;
	assert RAM(17682) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17682))))  severity failure;
	assert RAM(17683) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17683))))  severity failure;
	assert RAM(17684) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(17684))))  severity failure;
	assert RAM(17685) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(17685))))  severity failure;
	assert RAM(17686) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(17686))))  severity failure;
	assert RAM(17687) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(17687))))  severity failure;
	assert RAM(17688) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(17688))))  severity failure;
	assert RAM(17689) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17689))))  severity failure;
	assert RAM(17690) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(17690))))  severity failure;
	assert RAM(17691) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(17691))))  severity failure;
	assert RAM(17692) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(17692))))  severity failure;
	assert RAM(17693) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17693))))  severity failure;
	assert RAM(17694) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(17694))))  severity failure;
	assert RAM(17695) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(17695))))  severity failure;
	assert RAM(17696) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(17696))))  severity failure;
	assert RAM(17697) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17697))))  severity failure;
	assert RAM(17698) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17698))))  severity failure;
	assert RAM(17699) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(17699))))  severity failure;
	assert RAM(17700) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(17700))))  severity failure;
	assert RAM(17701) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(17701))))  severity failure;
	assert RAM(17702) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(17702))))  severity failure;
	assert RAM(17703) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17703))))  severity failure;
	assert RAM(17704) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(17704))))  severity failure;
	assert RAM(17705) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(17705))))  severity failure;
	assert RAM(17706) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(17706))))  severity failure;
	assert RAM(17707) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(17707))))  severity failure;
	assert RAM(17708) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(17708))))  severity failure;
	assert RAM(17709) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(17709))))  severity failure;
	assert RAM(17710) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17710))))  severity failure;
	assert RAM(17711) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(17711))))  severity failure;
	assert RAM(17712) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(17712))))  severity failure;
	assert RAM(17713) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17713))))  severity failure;
	assert RAM(17714) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(17714))))  severity failure;
	assert RAM(17715) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(17715))))  severity failure;
	assert RAM(17716) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(17716))))  severity failure;
	assert RAM(17717) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(17717))))  severity failure;
	assert RAM(17718) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(17718))))  severity failure;
	assert RAM(17719) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17719))))  severity failure;
	assert RAM(17720) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(17720))))  severity failure;
	assert RAM(17721) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17721))))  severity failure;
	assert RAM(17722) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(17722))))  severity failure;
	assert RAM(17723) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(17723))))  severity failure;
	assert RAM(17724) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(17724))))  severity failure;
	assert RAM(17725) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(17725))))  severity failure;
	assert RAM(17726) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17726))))  severity failure;
	assert RAM(17727) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(17727))))  severity failure;
	assert RAM(17728) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(17728))))  severity failure;
	assert RAM(17729) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(17729))))  severity failure;
	assert RAM(17730) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17730))))  severity failure;
	assert RAM(17731) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17731))))  severity failure;
	assert RAM(17732) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(17732))))  severity failure;
	assert RAM(17733) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(17733))))  severity failure;
	assert RAM(17734) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(17734))))  severity failure;
	assert RAM(17735) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(17735))))  severity failure;
	assert RAM(17736) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(17736))))  severity failure;
	assert RAM(17737) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17737))))  severity failure;
	assert RAM(17738) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17738))))  severity failure;
	assert RAM(17739) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(17739))))  severity failure;
	assert RAM(17740) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17740))))  severity failure;
	assert RAM(17741) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(17741))))  severity failure;
	assert RAM(17742) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(17742))))  severity failure;
	assert RAM(17743) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(17743))))  severity failure;
	assert RAM(17744) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(17744))))  severity failure;
	assert RAM(17745) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(17745))))  severity failure;
	assert RAM(17746) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17746))))  severity failure;
	assert RAM(17747) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(17747))))  severity failure;
	assert RAM(17748) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(17748))))  severity failure;
	assert RAM(17749) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17749))))  severity failure;
	assert RAM(17750) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(17750))))  severity failure;
	assert RAM(17751) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(17751))))  severity failure;
	assert RAM(17752) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(17752))))  severity failure;
	assert RAM(17753) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(17753))))  severity failure;
	assert RAM(17754) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(17754))))  severity failure;
	assert RAM(17755) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17755))))  severity failure;
	assert RAM(17756) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(17756))))  severity failure;
	assert RAM(17757) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(17757))))  severity failure;
	assert RAM(17758) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(17758))))  severity failure;
	assert RAM(17759) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17759))))  severity failure;
	assert RAM(17760) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(17760))))  severity failure;
	assert RAM(17761) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17761))))  severity failure;
	assert RAM(17762) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(17762))))  severity failure;
	assert RAM(17763) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(17763))))  severity failure;
	assert RAM(17764) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(17764))))  severity failure;
	assert RAM(17765) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(17765))))  severity failure;
	assert RAM(17766) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17766))))  severity failure;
	assert RAM(17767) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(17767))))  severity failure;
	assert RAM(17768) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(17768))))  severity failure;
	assert RAM(17769) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17769))))  severity failure;
	assert RAM(17770) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17770))))  severity failure;
	assert RAM(17771) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(17771))))  severity failure;
	assert RAM(17772) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17772))))  severity failure;
	assert RAM(17773) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(17773))))  severity failure;
	assert RAM(17774) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(17774))))  severity failure;
	assert RAM(17775) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17775))))  severity failure;
	assert RAM(17776) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(17776))))  severity failure;
	assert RAM(17777) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(17777))))  severity failure;
	assert RAM(17778) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(17778))))  severity failure;
	assert RAM(17779) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(17779))))  severity failure;
	assert RAM(17780) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(17780))))  severity failure;
	assert RAM(17781) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17781))))  severity failure;
	assert RAM(17782) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(17782))))  severity failure;
	assert RAM(17783) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(17783))))  severity failure;
	assert RAM(17784) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(17784))))  severity failure;
	assert RAM(17785) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(17785))))  severity failure;
	assert RAM(17786) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(17786))))  severity failure;
	assert RAM(17787) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(17787))))  severity failure;
	assert RAM(17788) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(17788))))  severity failure;
	assert RAM(17789) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(17789))))  severity failure;
	assert RAM(17790) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(17790))))  severity failure;
	assert RAM(17791) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(17791))))  severity failure;
	assert RAM(17792) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(17792))))  severity failure;
	assert RAM(17793) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(17793))))  severity failure;
	assert RAM(17794) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(17794))))  severity failure;
	assert RAM(17795) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(17795))))  severity failure;
	assert RAM(17796) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17796))))  severity failure;
	assert RAM(17797) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17797))))  severity failure;
	assert RAM(17798) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(17798))))  severity failure;
	assert RAM(17799) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(17799))))  severity failure;
	assert RAM(17800) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(17800))))  severity failure;
	assert RAM(17801) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(17801))))  severity failure;
	assert RAM(17802) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(17802))))  severity failure;
	assert RAM(17803) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(17803))))  severity failure;
	assert RAM(17804) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(17804))))  severity failure;
	assert RAM(17805) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(17805))))  severity failure;
	assert RAM(17806) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(17806))))  severity failure;
	assert RAM(17807) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(17807))))  severity failure;
	assert RAM(17808) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(17808))))  severity failure;
	assert RAM(17809) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(17809))))  severity failure;
	assert RAM(17810) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(17810))))  severity failure;
	assert RAM(17811) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17811))))  severity failure;
	assert RAM(17812) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17812))))  severity failure;
	assert RAM(17813) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17813))))  severity failure;
	assert RAM(17814) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17814))))  severity failure;
	assert RAM(17815) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(17815))))  severity failure;
	assert RAM(17816) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(17816))))  severity failure;
	assert RAM(17817) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(17817))))  severity failure;
	assert RAM(17818) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(17818))))  severity failure;
	assert RAM(17819) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17819))))  severity failure;
	assert RAM(17820) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(17820))))  severity failure;
	assert RAM(17821) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(17821))))  severity failure;
	assert RAM(17822) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(17822))))  severity failure;
	assert RAM(17823) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(17823))))  severity failure;
	assert RAM(17824) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(17824))))  severity failure;
	assert RAM(17825) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(17825))))  severity failure;
	assert RAM(17826) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17826))))  severity failure;
	assert RAM(17827) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(17827))))  severity failure;
	assert RAM(17828) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(17828))))  severity failure;
	assert RAM(17829) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17829))))  severity failure;
	assert RAM(17830) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(17830))))  severity failure;
	assert RAM(17831) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17831))))  severity failure;
	assert RAM(17832) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(17832))))  severity failure;
	assert RAM(17833) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17833))))  severity failure;
	assert RAM(17834) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(17834))))  severity failure;
	assert RAM(17835) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(17835))))  severity failure;
	assert RAM(17836) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(17836))))  severity failure;
	assert RAM(17837) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(17837))))  severity failure;
	assert RAM(17838) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(17838))))  severity failure;
	assert RAM(17839) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17839))))  severity failure;
	assert RAM(17840) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(17840))))  severity failure;
	assert RAM(17841) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17841))))  severity failure;
	assert RAM(17842) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(17842))))  severity failure;
	assert RAM(17843) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(17843))))  severity failure;
	assert RAM(17844) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(17844))))  severity failure;
	assert RAM(17845) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(17845))))  severity failure;
	assert RAM(17846) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(17846))))  severity failure;
	assert RAM(17847) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17847))))  severity failure;
	assert RAM(17848) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(17848))))  severity failure;
	assert RAM(17849) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17849))))  severity failure;
	assert RAM(17850) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(17850))))  severity failure;
	assert RAM(17851) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(17851))))  severity failure;
	assert RAM(17852) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(17852))))  severity failure;
	assert RAM(17853) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(17853))))  severity failure;
	assert RAM(17854) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(17854))))  severity failure;
	assert RAM(17855) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(17855))))  severity failure;
	assert RAM(17856) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(17856))))  severity failure;
	assert RAM(17857) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(17857))))  severity failure;
	assert RAM(17858) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(17858))))  severity failure;
	assert RAM(17859) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(17859))))  severity failure;
	assert RAM(17860) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(17860))))  severity failure;
	assert RAM(17861) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(17861))))  severity failure;
	assert RAM(17862) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(17862))))  severity failure;
	assert RAM(17863) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(17863))))  severity failure;
	assert RAM(17864) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(17864))))  severity failure;
	assert RAM(17865) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(17865))))  severity failure;
	assert RAM(17866) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(17866))))  severity failure;
	assert RAM(17867) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(17867))))  severity failure;
	assert RAM(17868) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(17868))))  severity failure;
	assert RAM(17869) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(17869))))  severity failure;
	assert RAM(17870) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(17870))))  severity failure;
	assert RAM(17871) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(17871))))  severity failure;
	assert RAM(17872) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(17872))))  severity failure;
	assert RAM(17873) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(17873))))  severity failure;
	assert RAM(17874) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(17874))))  severity failure;
	assert RAM(17875) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(17875))))  severity failure;
	assert RAM(17876) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(17876))))  severity failure;
	assert RAM(17877) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(17877))))  severity failure;
	assert RAM(17878) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(17878))))  severity failure;
	assert RAM(17879) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17879))))  severity failure;
	assert RAM(17880) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(17880))))  severity failure;
	assert RAM(17881) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(17881))))  severity failure;
	assert RAM(17882) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(17882))))  severity failure;
	assert RAM(17883) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(17883))))  severity failure;
	assert RAM(17884) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(17884))))  severity failure;
	assert RAM(17885) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(17885))))  severity failure;
	assert RAM(17886) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(17886))))  severity failure;
	assert RAM(17887) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(17887))))  severity failure;
	assert RAM(17888) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(17888))))  severity failure;
	assert RAM(17889) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(17889))))  severity failure;
	assert RAM(17890) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(17890))))  severity failure;
	assert RAM(17891) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(17891))))  severity failure;
	assert RAM(17892) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(17892))))  severity failure;
	assert RAM(17893) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(17893))))  severity failure;
	assert RAM(17894) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(17894))))  severity failure;
	assert RAM(17895) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(17895))))  severity failure;
	assert RAM(17896) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(17896))))  severity failure;
	assert RAM(17897) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(17897))))  severity failure;
	assert RAM(17898) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(17898))))  severity failure;
	assert RAM(17899) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(17899))))  severity failure;
	assert RAM(17900) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(17900))))  severity failure;
	assert RAM(17901) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(17901))))  severity failure;
	assert RAM(17902) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(17902))))  severity failure;
	assert RAM(17903) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(17903))))  severity failure;
	assert RAM(17904) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(17904))))  severity failure;
	assert RAM(17905) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(17905))))  severity failure;
	assert RAM(17906) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(17906))))  severity failure;
	assert RAM(17907) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(17907))))  severity failure;
	assert RAM(17908) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(17908))))  severity failure;
	assert RAM(17909) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(17909))))  severity failure;
	assert RAM(17910) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(17910))))  severity failure;
	assert RAM(17911) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(17911))))  severity failure;
	assert RAM(17912) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(17912))))  severity failure;
	assert RAM(17913) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(17913))))  severity failure;
	assert RAM(17914) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(17914))))  severity failure;
	assert RAM(17915) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(17915))))  severity failure;
	assert RAM(17916) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(17916))))  severity failure;
	assert RAM(17917) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(17917))))  severity failure;
	assert RAM(17918) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(17918))))  severity failure;
	assert RAM(17919) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(17919))))  severity failure;
	assert RAM(17920) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(17920))))  severity failure;
	assert RAM(17921) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17921))))  severity failure;
	assert RAM(17922) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(17922))))  severity failure;
	assert RAM(17923) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(17923))))  severity failure;
	assert RAM(17924) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(17924))))  severity failure;
	assert RAM(17925) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(17925))))  severity failure;
	assert RAM(17926) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(17926))))  severity failure;
	assert RAM(17927) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(17927))))  severity failure;
	assert RAM(17928) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(17928))))  severity failure;
	assert RAM(17929) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(17929))))  severity failure;
	assert RAM(17930) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(17930))))  severity failure;
	assert RAM(17931) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17931))))  severity failure;
	assert RAM(17932) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(17932))))  severity failure;
	assert RAM(17933) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(17933))))  severity failure;
	assert RAM(17934) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17934))))  severity failure;
	assert RAM(17935) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(17935))))  severity failure;
	assert RAM(17936) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(17936))))  severity failure;
	assert RAM(17937) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(17937))))  severity failure;
	assert RAM(17938) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(17938))))  severity failure;
	assert RAM(17939) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(17939))))  severity failure;
	assert RAM(17940) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(17940))))  severity failure;
	assert RAM(17941) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(17941))))  severity failure;
	assert RAM(17942) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(17942))))  severity failure;
	assert RAM(17943) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(17943))))  severity failure;
	assert RAM(17944) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(17944))))  severity failure;
	assert RAM(17945) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(17945))))  severity failure;
	assert RAM(17946) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(17946))))  severity failure;
	assert RAM(17947) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(17947))))  severity failure;
	assert RAM(17948) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(17948))))  severity failure;
	assert RAM(17949) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(17949))))  severity failure;
	assert RAM(17950) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(17950))))  severity failure;
	assert RAM(17951) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(17951))))  severity failure;
	assert RAM(17952) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(17952))))  severity failure;
	assert RAM(17953) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(17953))))  severity failure;
	assert RAM(17954) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(17954))))  severity failure;
	assert RAM(17955) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(17955))))  severity failure;
	assert RAM(17956) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(17956))))  severity failure;
	assert RAM(17957) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(17957))))  severity failure;
	assert RAM(17958) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(17958))))  severity failure;
	assert RAM(17959) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(17959))))  severity failure;
	assert RAM(17960) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(17960))))  severity failure;
	assert RAM(17961) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(17961))))  severity failure;
	assert RAM(17962) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(17962))))  severity failure;
	assert RAM(17963) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(17963))))  severity failure;
	assert RAM(17964) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(17964))))  severity failure;
	assert RAM(17965) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(17965))))  severity failure;
	assert RAM(17966) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(17966))))  severity failure;
	assert RAM(17967) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(17967))))  severity failure;
	assert RAM(17968) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(17968))))  severity failure;
	assert RAM(17969) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(17969))))  severity failure;
	assert RAM(17970) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(17970))))  severity failure;
	assert RAM(17971) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(17971))))  severity failure;
	assert RAM(17972) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(17972))))  severity failure;
	assert RAM(17973) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(17973))))  severity failure;
	assert RAM(17974) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(17974))))  severity failure;
	assert RAM(17975) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(17975))))  severity failure;
	assert RAM(17976) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(17976))))  severity failure;
	assert RAM(17977) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(17977))))  severity failure;
	assert RAM(17978) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(17978))))  severity failure;
	assert RAM(17979) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(17979))))  severity failure;
	assert RAM(17980) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(17980))))  severity failure;
	assert RAM(17981) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(17981))))  severity failure;
	assert RAM(17982) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(17982))))  severity failure;
	assert RAM(17983) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(17983))))  severity failure;
	assert RAM(17984) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(17984))))  severity failure;
	assert RAM(17985) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(17985))))  severity failure;
	assert RAM(17986) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(17986))))  severity failure;
	assert RAM(17987) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(17987))))  severity failure;
	assert RAM(17988) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(17988))))  severity failure;
	assert RAM(17989) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(17989))))  severity failure;
	assert RAM(17990) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(17990))))  severity failure;
	assert RAM(17991) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(17991))))  severity failure;
	assert RAM(17992) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(17992))))  severity failure;
	assert RAM(17993) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(17993))))  severity failure;
	assert RAM(17994) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(17994))))  severity failure;
	assert RAM(17995) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(17995))))  severity failure;
	assert RAM(17996) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(17996))))  severity failure;
	assert RAM(17997) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(17997))))  severity failure;
	assert RAM(17998) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(17998))))  severity failure;
	assert RAM(17999) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(17999))))  severity failure;
	assert RAM(18000) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(18000))))  severity failure;
	assert RAM(18001) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18001))))  severity failure;
	assert RAM(18002) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18002))))  severity failure;
	assert RAM(18003) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18003))))  severity failure;
	assert RAM(18004) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18004))))  severity failure;
	assert RAM(18005) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(18005))))  severity failure;
	assert RAM(18006) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(18006))))  severity failure;
	assert RAM(18007) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18007))))  severity failure;
	assert RAM(18008) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(18008))))  severity failure;
	assert RAM(18009) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(18009))))  severity failure;
	assert RAM(18010) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(18010))))  severity failure;
	assert RAM(18011) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18011))))  severity failure;
	assert RAM(18012) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18012))))  severity failure;
	assert RAM(18013) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(18013))))  severity failure;
	assert RAM(18014) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(18014))))  severity failure;
	assert RAM(18015) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(18015))))  severity failure;
	assert RAM(18016) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(18016))))  severity failure;
	assert RAM(18017) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(18017))))  severity failure;
	assert RAM(18018) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(18018))))  severity failure;
	assert RAM(18019) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(18019))))  severity failure;
	assert RAM(18020) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18020))))  severity failure;
	assert RAM(18021) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(18021))))  severity failure;
	assert RAM(18022) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(18022))))  severity failure;
	assert RAM(18023) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18023))))  severity failure;
	assert RAM(18024) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(18024))))  severity failure;
	assert RAM(18025) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18025))))  severity failure;
	assert RAM(18026) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(18026))))  severity failure;
	assert RAM(18027) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(18027))))  severity failure;
	assert RAM(18028) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18028))))  severity failure;
	assert RAM(18029) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(18029))))  severity failure;
	assert RAM(18030) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(18030))))  severity failure;
	assert RAM(18031) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(18031))))  severity failure;
	assert RAM(18032) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18032))))  severity failure;
	assert RAM(18033) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(18033))))  severity failure;
	assert RAM(18034) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(18034))))  severity failure;
	assert RAM(18035) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(18035))))  severity failure;
	assert RAM(18036) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18036))))  severity failure;
	assert RAM(18037) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18037))))  severity failure;
	assert RAM(18038) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(18038))))  severity failure;
	assert RAM(18039) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(18039))))  severity failure;
	assert RAM(18040) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18040))))  severity failure;
	assert RAM(18041) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(18041))))  severity failure;
	assert RAM(18042) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(18042))))  severity failure;
	assert RAM(18043) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(18043))))  severity failure;
	assert RAM(18044) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(18044))))  severity failure;
	assert RAM(18045) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(18045))))  severity failure;
	assert RAM(18046) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(18046))))  severity failure;
	assert RAM(18047) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(18047))))  severity failure;
	assert RAM(18048) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(18048))))  severity failure;
	assert RAM(18049) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(18049))))  severity failure;
	assert RAM(18050) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(18050))))  severity failure;
	assert RAM(18051) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(18051))))  severity failure;
	assert RAM(18052) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(18052))))  severity failure;
	assert RAM(18053) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(18053))))  severity failure;
	assert RAM(18054) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18054))))  severity failure;
	assert RAM(18055) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18055))))  severity failure;
	assert RAM(18056) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(18056))))  severity failure;
	assert RAM(18057) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18057))))  severity failure;
	assert RAM(18058) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(18058))))  severity failure;
	assert RAM(18059) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18059))))  severity failure;
	assert RAM(18060) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(18060))))  severity failure;
	assert RAM(18061) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(18061))))  severity failure;
	assert RAM(18062) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(18062))))  severity failure;
	assert RAM(18063) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(18063))))  severity failure;
	assert RAM(18064) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(18064))))  severity failure;
	assert RAM(18065) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18065))))  severity failure;
	assert RAM(18066) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(18066))))  severity failure;
	assert RAM(18067) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18067))))  severity failure;
	assert RAM(18068) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(18068))))  severity failure;
	assert RAM(18069) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(18069))))  severity failure;
	assert RAM(18070) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(18070))))  severity failure;
	assert RAM(18071) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(18071))))  severity failure;
	assert RAM(18072) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18072))))  severity failure;
	assert RAM(18073) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(18073))))  severity failure;
	assert RAM(18074) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(18074))))  severity failure;
	assert RAM(18075) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(18075))))  severity failure;
	assert RAM(18076) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(18076))))  severity failure;
	assert RAM(18077) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(18077))))  severity failure;
	assert RAM(18078) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(18078))))  severity failure;
	assert RAM(18079) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(18079))))  severity failure;
	assert RAM(18080) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18080))))  severity failure;
	assert RAM(18081) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(18081))))  severity failure;
	assert RAM(18082) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(18082))))  severity failure;
	assert RAM(18083) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(18083))))  severity failure;
	assert RAM(18084) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18084))))  severity failure;
	assert RAM(18085) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(18085))))  severity failure;
	assert RAM(18086) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18086))))  severity failure;
	assert RAM(18087) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18087))))  severity failure;
	assert RAM(18088) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18088))))  severity failure;
	assert RAM(18089) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(18089))))  severity failure;
	assert RAM(18090) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(18090))))  severity failure;
	assert RAM(18091) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(18091))))  severity failure;
	assert RAM(18092) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(18092))))  severity failure;
	assert RAM(18093) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18093))))  severity failure;
	assert RAM(18094) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(18094))))  severity failure;
	assert RAM(18095) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(18095))))  severity failure;
	assert RAM(18096) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(18096))))  severity failure;
	assert RAM(18097) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(18097))))  severity failure;
	assert RAM(18098) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(18098))))  severity failure;
	assert RAM(18099) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(18099))))  severity failure;
	assert RAM(18100) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(18100))))  severity failure;
	assert RAM(18101) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(18101))))  severity failure;
	assert RAM(18102) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(18102))))  severity failure;
	assert RAM(18103) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(18103))))  severity failure;
	assert RAM(18104) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(18104))))  severity failure;
	assert RAM(18105) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(18105))))  severity failure;
	assert RAM(18106) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(18106))))  severity failure;
	assert RAM(18107) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18107))))  severity failure;
	assert RAM(18108) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18108))))  severity failure;
	assert RAM(18109) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18109))))  severity failure;
	assert RAM(18110) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(18110))))  severity failure;
	assert RAM(18111) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(18111))))  severity failure;
	assert RAM(18112) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(18112))))  severity failure;
	assert RAM(18113) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(18113))))  severity failure;
	assert RAM(18114) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(18114))))  severity failure;
	assert RAM(18115) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(18115))))  severity failure;
	assert RAM(18116) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(18116))))  severity failure;
	assert RAM(18117) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18117))))  severity failure;
	assert RAM(18118) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18118))))  severity failure;
	assert RAM(18119) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18119))))  severity failure;
	assert RAM(18120) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(18120))))  severity failure;
	assert RAM(18121) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(18121))))  severity failure;
	assert RAM(18122) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(18122))))  severity failure;
	assert RAM(18123) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(18123))))  severity failure;
	assert RAM(18124) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(18124))))  severity failure;
	assert RAM(18125) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18125))))  severity failure;
	assert RAM(18126) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(18126))))  severity failure;
	assert RAM(18127) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(18127))))  severity failure;
	assert RAM(18128) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18128))))  severity failure;
	assert RAM(18129) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(18129))))  severity failure;
	assert RAM(18130) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18130))))  severity failure;
	assert RAM(18131) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(18131))))  severity failure;
	assert RAM(18132) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(18132))))  severity failure;
	assert RAM(18133) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(18133))))  severity failure;
	assert RAM(18134) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(18134))))  severity failure;
	assert RAM(18135) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18135))))  severity failure;
	assert RAM(18136) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(18136))))  severity failure;
	assert RAM(18137) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(18137))))  severity failure;
	assert RAM(18138) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18138))))  severity failure;
	assert RAM(18139) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(18139))))  severity failure;
	assert RAM(18140) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(18140))))  severity failure;
	assert RAM(18141) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(18141))))  severity failure;
	assert RAM(18142) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(18142))))  severity failure;
	assert RAM(18143) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(18143))))  severity failure;
	assert RAM(18144) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(18144))))  severity failure;
	assert RAM(18145) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(18145))))  severity failure;
	assert RAM(18146) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(18146))))  severity failure;
	assert RAM(18147) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(18147))))  severity failure;
	assert RAM(18148) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18148))))  severity failure;
	assert RAM(18149) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(18149))))  severity failure;
	assert RAM(18150) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18150))))  severity failure;
	assert RAM(18151) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18151))))  severity failure;
	assert RAM(18152) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18152))))  severity failure;
	assert RAM(18153) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(18153))))  severity failure;
	assert RAM(18154) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(18154))))  severity failure;
	assert RAM(18155) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(18155))))  severity failure;
	assert RAM(18156) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(18156))))  severity failure;
	assert RAM(18157) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(18157))))  severity failure;
	assert RAM(18158) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(18158))))  severity failure;
	assert RAM(18159) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18159))))  severity failure;
	assert RAM(18160) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(18160))))  severity failure;
	assert RAM(18161) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(18161))))  severity failure;
	assert RAM(18162) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(18162))))  severity failure;
	assert RAM(18163) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18163))))  severity failure;
	assert RAM(18164) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18164))))  severity failure;
	assert RAM(18165) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(18165))))  severity failure;
	assert RAM(18166) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(18166))))  severity failure;
	assert RAM(18167) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18167))))  severity failure;
	assert RAM(18168) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18168))))  severity failure;
	assert RAM(18169) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(18169))))  severity failure;
	assert RAM(18170) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18170))))  severity failure;
	assert RAM(18171) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(18171))))  severity failure;
	assert RAM(18172) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18172))))  severity failure;
	assert RAM(18173) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18173))))  severity failure;
	assert RAM(18174) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(18174))))  severity failure;
	assert RAM(18175) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18175))))  severity failure;
	assert RAM(18176) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(18176))))  severity failure;
	assert RAM(18177) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(18177))))  severity failure;
	assert RAM(18178) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(18178))))  severity failure;
	assert RAM(18179) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(18179))))  severity failure;
	assert RAM(18180) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(18180))))  severity failure;
	assert RAM(18181) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(18181))))  severity failure;
	assert RAM(18182) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18182))))  severity failure;
	assert RAM(18183) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(18183))))  severity failure;
	assert RAM(18184) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(18184))))  severity failure;
	assert RAM(18185) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(18185))))  severity failure;
	assert RAM(18186) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(18186))))  severity failure;
	assert RAM(18187) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(18187))))  severity failure;
	assert RAM(18188) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(18188))))  severity failure;
	assert RAM(18189) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18189))))  severity failure;
	assert RAM(18190) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(18190))))  severity failure;
	assert RAM(18191) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(18191))))  severity failure;
	assert RAM(18192) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(18192))))  severity failure;
	assert RAM(18193) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(18193))))  severity failure;
	assert RAM(18194) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(18194))))  severity failure;
	assert RAM(18195) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(18195))))  severity failure;
	assert RAM(18196) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(18196))))  severity failure;
	assert RAM(18197) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18197))))  severity failure;
	assert RAM(18198) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(18198))))  severity failure;
	assert RAM(18199) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18199))))  severity failure;
	assert RAM(18200) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(18200))))  severity failure;
	assert RAM(18201) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(18201))))  severity failure;
	assert RAM(18202) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18202))))  severity failure;
	assert RAM(18203) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(18203))))  severity failure;
	assert RAM(18204) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(18204))))  severity failure;
	assert RAM(18205) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(18205))))  severity failure;
	assert RAM(18206) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(18206))))  severity failure;
	assert RAM(18207) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18207))))  severity failure;
	assert RAM(18208) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(18208))))  severity failure;
	assert RAM(18209) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18209))))  severity failure;
	assert RAM(18210) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(18210))))  severity failure;
	assert RAM(18211) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(18211))))  severity failure;
	assert RAM(18212) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(18212))))  severity failure;
	assert RAM(18213) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(18213))))  severity failure;
	assert RAM(18214) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18214))))  severity failure;
	assert RAM(18215) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(18215))))  severity failure;
	assert RAM(18216) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(18216))))  severity failure;
	assert RAM(18217) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18217))))  severity failure;
	assert RAM(18218) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(18218))))  severity failure;
	assert RAM(18219) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(18219))))  severity failure;
	assert RAM(18220) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(18220))))  severity failure;
	assert RAM(18221) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18221))))  severity failure;
	assert RAM(18222) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(18222))))  severity failure;
	assert RAM(18223) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(18223))))  severity failure;
	assert RAM(18224) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(18224))))  severity failure;
	assert RAM(18225) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18225))))  severity failure;
	assert RAM(18226) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18226))))  severity failure;
	assert RAM(18227) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18227))))  severity failure;
	assert RAM(18228) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18228))))  severity failure;
	assert RAM(18229) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(18229))))  severity failure;
	assert RAM(18230) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18230))))  severity failure;
	assert RAM(18231) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(18231))))  severity failure;
	assert RAM(18232) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(18232))))  severity failure;
	assert RAM(18233) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(18233))))  severity failure;
	assert RAM(18234) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(18234))))  severity failure;
	assert RAM(18235) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(18235))))  severity failure;
	assert RAM(18236) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(18236))))  severity failure;
	assert RAM(18237) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(18237))))  severity failure;
	assert RAM(18238) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(18238))))  severity failure;
	assert RAM(18239) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18239))))  severity failure;
	assert RAM(18240) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(18240))))  severity failure;
	assert RAM(18241) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(18241))))  severity failure;
	assert RAM(18242) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(18242))))  severity failure;
	assert RAM(18243) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(18243))))  severity failure;
	assert RAM(18244) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(18244))))  severity failure;
	assert RAM(18245) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(18245))))  severity failure;
	assert RAM(18246) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(18246))))  severity failure;
	assert RAM(18247) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18247))))  severity failure;
	assert RAM(18248) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18248))))  severity failure;
	assert RAM(18249) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(18249))))  severity failure;
	assert RAM(18250) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(18250))))  severity failure;
	assert RAM(18251) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(18251))))  severity failure;
	assert RAM(18252) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(18252))))  severity failure;
	assert RAM(18253) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(18253))))  severity failure;
	assert RAM(18254) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(18254))))  severity failure;
	assert RAM(18255) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(18255))))  severity failure;
	assert RAM(18256) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18256))))  severity failure;
	assert RAM(18257) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18257))))  severity failure;
	assert RAM(18258) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(18258))))  severity failure;
	assert RAM(18259) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(18259))))  severity failure;
	assert RAM(18260) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(18260))))  severity failure;
	assert RAM(18261) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(18261))))  severity failure;
	assert RAM(18262) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(18262))))  severity failure;
	assert RAM(18263) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18263))))  severity failure;
	assert RAM(18264) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(18264))))  severity failure;
	assert RAM(18265) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(18265))))  severity failure;
	assert RAM(18266) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(18266))))  severity failure;
	assert RAM(18267) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(18267))))  severity failure;
	assert RAM(18268) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18268))))  severity failure;
	assert RAM(18269) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18269))))  severity failure;
	assert RAM(18270) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(18270))))  severity failure;
	assert RAM(18271) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(18271))))  severity failure;
	assert RAM(18272) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(18272))))  severity failure;
	assert RAM(18273) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(18273))))  severity failure;
	assert RAM(18274) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18274))))  severity failure;
	assert RAM(18275) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(18275))))  severity failure;
	assert RAM(18276) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18276))))  severity failure;
	assert RAM(18277) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18277))))  severity failure;
	assert RAM(18278) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(18278))))  severity failure;
	assert RAM(18279) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(18279))))  severity failure;
	assert RAM(18280) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(18280))))  severity failure;
	assert RAM(18281) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(18281))))  severity failure;
	assert RAM(18282) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(18282))))  severity failure;
	assert RAM(18283) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(18283))))  severity failure;
	assert RAM(18284) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(18284))))  severity failure;
	assert RAM(18285) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18285))))  severity failure;
	assert RAM(18286) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(18286))))  severity failure;
	assert RAM(18287) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(18287))))  severity failure;
	assert RAM(18288) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(18288))))  severity failure;
	assert RAM(18289) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(18289))))  severity failure;
	assert RAM(18290) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18290))))  severity failure;
	assert RAM(18291) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18291))))  severity failure;
	assert RAM(18292) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(18292))))  severity failure;
	assert RAM(18293) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(18293))))  severity failure;
	assert RAM(18294) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(18294))))  severity failure;
	assert RAM(18295) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(18295))))  severity failure;
	assert RAM(18296) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18296))))  severity failure;
	assert RAM(18297) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(18297))))  severity failure;
	assert RAM(18298) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18298))))  severity failure;
	assert RAM(18299) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(18299))))  severity failure;
	assert RAM(18300) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(18300))))  severity failure;
	assert RAM(18301) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(18301))))  severity failure;
	assert RAM(18302) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(18302))))  severity failure;
	assert RAM(18303) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(18303))))  severity failure;
	assert RAM(18304) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(18304))))  severity failure;
	assert RAM(18305) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(18305))))  severity failure;
	assert RAM(18306) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(18306))))  severity failure;
	assert RAM(18307) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(18307))))  severity failure;
	assert RAM(18308) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(18308))))  severity failure;
	assert RAM(18309) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18309))))  severity failure;
	assert RAM(18310) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(18310))))  severity failure;
	assert RAM(18311) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(18311))))  severity failure;
	assert RAM(18312) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18312))))  severity failure;
	assert RAM(18313) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(18313))))  severity failure;
	assert RAM(18314) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(18314))))  severity failure;
	assert RAM(18315) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(18315))))  severity failure;
	assert RAM(18316) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(18316))))  severity failure;
	assert RAM(18317) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(18317))))  severity failure;
	assert RAM(18318) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18318))))  severity failure;
	assert RAM(18319) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(18319))))  severity failure;
	assert RAM(18320) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18320))))  severity failure;
	assert RAM(18321) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(18321))))  severity failure;
	assert RAM(18322) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18322))))  severity failure;
	assert RAM(18323) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(18323))))  severity failure;
	assert RAM(18324) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(18324))))  severity failure;
	assert RAM(18325) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(18325))))  severity failure;
	assert RAM(18326) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18326))))  severity failure;
	assert RAM(18327) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(18327))))  severity failure;
	assert RAM(18328) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18328))))  severity failure;
	assert RAM(18329) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18329))))  severity failure;
	assert RAM(18330) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(18330))))  severity failure;
	assert RAM(18331) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18331))))  severity failure;
	assert RAM(18332) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18332))))  severity failure;
	assert RAM(18333) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18333))))  severity failure;
	assert RAM(18334) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18334))))  severity failure;
	assert RAM(18335) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(18335))))  severity failure;
	assert RAM(18336) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(18336))))  severity failure;
	assert RAM(18337) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(18337))))  severity failure;
	assert RAM(18338) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18338))))  severity failure;
	assert RAM(18339) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18339))))  severity failure;
	assert RAM(18340) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18340))))  severity failure;
	assert RAM(18341) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(18341))))  severity failure;
	assert RAM(18342) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18342))))  severity failure;
	assert RAM(18343) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(18343))))  severity failure;
	assert RAM(18344) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18344))))  severity failure;
	assert RAM(18345) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18345))))  severity failure;
	assert RAM(18346) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(18346))))  severity failure;
	assert RAM(18347) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(18347))))  severity failure;
	assert RAM(18348) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(18348))))  severity failure;
	assert RAM(18349) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18349))))  severity failure;
	assert RAM(18350) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(18350))))  severity failure;
	assert RAM(18351) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(18351))))  severity failure;
	assert RAM(18352) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(18352))))  severity failure;
	assert RAM(18353) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18353))))  severity failure;
	assert RAM(18354) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18354))))  severity failure;
	assert RAM(18355) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(18355))))  severity failure;
	assert RAM(18356) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(18356))))  severity failure;
	assert RAM(18357) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(18357))))  severity failure;
	assert RAM(18358) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(18358))))  severity failure;
	assert RAM(18359) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18359))))  severity failure;
	assert RAM(18360) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18360))))  severity failure;
	assert RAM(18361) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18361))))  severity failure;
	assert RAM(18362) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(18362))))  severity failure;
	assert RAM(18363) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(18363))))  severity failure;
	assert RAM(18364) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(18364))))  severity failure;
	assert RAM(18365) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(18365))))  severity failure;
	assert RAM(18366) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18366))))  severity failure;
	assert RAM(18367) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(18367))))  severity failure;
	assert RAM(18368) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18368))))  severity failure;
	assert RAM(18369) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(18369))))  severity failure;
	assert RAM(18370) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(18370))))  severity failure;
	assert RAM(18371) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(18371))))  severity failure;
	assert RAM(18372) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(18372))))  severity failure;
	assert RAM(18373) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(18373))))  severity failure;
	assert RAM(18374) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(18374))))  severity failure;
	assert RAM(18375) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(18375))))  severity failure;
	assert RAM(18376) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(18376))))  severity failure;
	assert RAM(18377) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(18377))))  severity failure;
	assert RAM(18378) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(18378))))  severity failure;
	assert RAM(18379) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(18379))))  severity failure;
	assert RAM(18380) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(18380))))  severity failure;
	assert RAM(18381) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(18381))))  severity failure;
	assert RAM(18382) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18382))))  severity failure;
	assert RAM(18383) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18383))))  severity failure;
	assert RAM(18384) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(18384))))  severity failure;
	assert RAM(18385) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(18385))))  severity failure;
	assert RAM(18386) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(18386))))  severity failure;
	assert RAM(18387) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(18387))))  severity failure;
	assert RAM(18388) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(18388))))  severity failure;
	assert RAM(18389) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(18389))))  severity failure;
	assert RAM(18390) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18390))))  severity failure;
	assert RAM(18391) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(18391))))  severity failure;
	assert RAM(18392) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(18392))))  severity failure;
	assert RAM(18393) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(18393))))  severity failure;
	assert RAM(18394) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18394))))  severity failure;
	assert RAM(18395) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18395))))  severity failure;
	assert RAM(18396) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(18396))))  severity failure;
	assert RAM(18397) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(18397))))  severity failure;
	assert RAM(18398) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(18398))))  severity failure;
	assert RAM(18399) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(18399))))  severity failure;
	assert RAM(18400) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(18400))))  severity failure;
	assert RAM(18401) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18401))))  severity failure;
	assert RAM(18402) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(18402))))  severity failure;
	assert RAM(18403) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(18403))))  severity failure;
	assert RAM(18404) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(18404))))  severity failure;
	assert RAM(18405) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(18405))))  severity failure;
	assert RAM(18406) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(18406))))  severity failure;
	assert RAM(18407) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(18407))))  severity failure;
	assert RAM(18408) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18408))))  severity failure;
	assert RAM(18409) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(18409))))  severity failure;
	assert RAM(18410) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(18410))))  severity failure;
	assert RAM(18411) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18411))))  severity failure;
	assert RAM(18412) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(18412))))  severity failure;
	assert RAM(18413) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(18413))))  severity failure;
	assert RAM(18414) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(18414))))  severity failure;
	assert RAM(18415) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(18415))))  severity failure;
	assert RAM(18416) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(18416))))  severity failure;
	assert RAM(18417) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(18417))))  severity failure;
	assert RAM(18418) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(18418))))  severity failure;
	assert RAM(18419) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(18419))))  severity failure;
	assert RAM(18420) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(18420))))  severity failure;
	assert RAM(18421) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(18421))))  severity failure;
	assert RAM(18422) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18422))))  severity failure;
	assert RAM(18423) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(18423))))  severity failure;
	assert RAM(18424) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(18424))))  severity failure;
	assert RAM(18425) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(18425))))  severity failure;
	assert RAM(18426) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(18426))))  severity failure;
	assert RAM(18427) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18427))))  severity failure;
	assert RAM(18428) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18428))))  severity failure;
	assert RAM(18429) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(18429))))  severity failure;
	assert RAM(18430) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(18430))))  severity failure;
	assert RAM(18431) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(18431))))  severity failure;
	assert RAM(18432) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(18432))))  severity failure;
	assert RAM(18433) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18433))))  severity failure;
	assert RAM(18434) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(18434))))  severity failure;
	assert RAM(18435) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(18435))))  severity failure;
	assert RAM(18436) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(18436))))  severity failure;
	assert RAM(18437) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(18437))))  severity failure;
	assert RAM(18438) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(18438))))  severity failure;
	assert RAM(18439) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(18439))))  severity failure;
	assert RAM(18440) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18440))))  severity failure;
	assert RAM(18441) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(18441))))  severity failure;
	assert RAM(18442) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(18442))))  severity failure;
	assert RAM(18443) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18443))))  severity failure;
	assert RAM(18444) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(18444))))  severity failure;
	assert RAM(18445) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(18445))))  severity failure;
	assert RAM(18446) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(18446))))  severity failure;
	assert RAM(18447) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(18447))))  severity failure;
	assert RAM(18448) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18448))))  severity failure;
	assert RAM(18449) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18449))))  severity failure;
	assert RAM(18450) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(18450))))  severity failure;
	assert RAM(18451) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(18451))))  severity failure;
	assert RAM(18452) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(18452))))  severity failure;
	assert RAM(18453) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(18453))))  severity failure;
	assert RAM(18454) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18454))))  severity failure;
	assert RAM(18455) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18455))))  severity failure;
	assert RAM(18456) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(18456))))  severity failure;
	assert RAM(18457) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(18457))))  severity failure;
	assert RAM(18458) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18458))))  severity failure;
	assert RAM(18459) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(18459))))  severity failure;
	assert RAM(18460) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(18460))))  severity failure;
	assert RAM(18461) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(18461))))  severity failure;
	assert RAM(18462) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(18462))))  severity failure;
	assert RAM(18463) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(18463))))  severity failure;
	assert RAM(18464) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18464))))  severity failure;
	assert RAM(18465) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(18465))))  severity failure;
	assert RAM(18466) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18466))))  severity failure;
	assert RAM(18467) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(18467))))  severity failure;
	assert RAM(18468) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(18468))))  severity failure;
	assert RAM(18469) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(18469))))  severity failure;
	assert RAM(18470) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18470))))  severity failure;
	assert RAM(18471) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(18471))))  severity failure;
	assert RAM(18472) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(18472))))  severity failure;
	assert RAM(18473) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18473))))  severity failure;
	assert RAM(18474) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(18474))))  severity failure;
	assert RAM(18475) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(18475))))  severity failure;
	assert RAM(18476) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(18476))))  severity failure;
	assert RAM(18477) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(18477))))  severity failure;
	assert RAM(18478) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(18478))))  severity failure;
	assert RAM(18479) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(18479))))  severity failure;
	assert RAM(18480) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18480))))  severity failure;
	assert RAM(18481) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(18481))))  severity failure;
	assert RAM(18482) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18482))))  severity failure;
	assert RAM(18483) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(18483))))  severity failure;
	assert RAM(18484) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18484))))  severity failure;
	assert RAM(18485) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(18485))))  severity failure;
	assert RAM(18486) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(18486))))  severity failure;
	assert RAM(18487) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(18487))))  severity failure;
	assert RAM(18488) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(18488))))  severity failure;
	assert RAM(18489) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18489))))  severity failure;
	assert RAM(18490) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(18490))))  severity failure;
	assert RAM(18491) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18491))))  severity failure;
	assert RAM(18492) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(18492))))  severity failure;
	assert RAM(18493) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18493))))  severity failure;
	assert RAM(18494) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(18494))))  severity failure;
	assert RAM(18495) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(18495))))  severity failure;
	assert RAM(18496) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(18496))))  severity failure;
	assert RAM(18497) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18497))))  severity failure;
	assert RAM(18498) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(18498))))  severity failure;
	assert RAM(18499) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(18499))))  severity failure;
	assert RAM(18500) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(18500))))  severity failure;
	assert RAM(18501) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(18501))))  severity failure;
	assert RAM(18502) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18502))))  severity failure;
	assert RAM(18503) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18503))))  severity failure;
	assert RAM(18504) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(18504))))  severity failure;
	assert RAM(18505) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(18505))))  severity failure;
	assert RAM(18506) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(18506))))  severity failure;
	assert RAM(18507) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(18507))))  severity failure;
	assert RAM(18508) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(18508))))  severity failure;
	assert RAM(18509) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(18509))))  severity failure;
	assert RAM(18510) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(18510))))  severity failure;
	assert RAM(18511) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(18511))))  severity failure;
	assert RAM(18512) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(18512))))  severity failure;
	assert RAM(18513) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18513))))  severity failure;
	assert RAM(18514) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(18514))))  severity failure;
	assert RAM(18515) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(18515))))  severity failure;
	assert RAM(18516) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(18516))))  severity failure;
	assert RAM(18517) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(18517))))  severity failure;
	assert RAM(18518) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(18518))))  severity failure;
	assert RAM(18519) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18519))))  severity failure;
	assert RAM(18520) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(18520))))  severity failure;
	assert RAM(18521) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18521))))  severity failure;
	assert RAM(18522) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(18522))))  severity failure;
	assert RAM(18523) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18523))))  severity failure;
	assert RAM(18524) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(18524))))  severity failure;
	assert RAM(18525) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(18525))))  severity failure;
	assert RAM(18526) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(18526))))  severity failure;
	assert RAM(18527) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(18527))))  severity failure;
	assert RAM(18528) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(18528))))  severity failure;
	assert RAM(18529) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(18529))))  severity failure;
	assert RAM(18530) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(18530))))  severity failure;
	assert RAM(18531) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(18531))))  severity failure;
	assert RAM(18532) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18532))))  severity failure;
	assert RAM(18533) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(18533))))  severity failure;
	assert RAM(18534) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(18534))))  severity failure;
	assert RAM(18535) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(18535))))  severity failure;
	assert RAM(18536) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(18536))))  severity failure;
	assert RAM(18537) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18537))))  severity failure;
	assert RAM(18538) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18538))))  severity failure;
	assert RAM(18539) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18539))))  severity failure;
	assert RAM(18540) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18540))))  severity failure;
	assert RAM(18541) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18541))))  severity failure;
	assert RAM(18542) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(18542))))  severity failure;
	assert RAM(18543) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(18543))))  severity failure;
	assert RAM(18544) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(18544))))  severity failure;
	assert RAM(18545) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18545))))  severity failure;
	assert RAM(18546) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(18546))))  severity failure;
	assert RAM(18547) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(18547))))  severity failure;
	assert RAM(18548) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18548))))  severity failure;
	assert RAM(18549) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18549))))  severity failure;
	assert RAM(18550) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(18550))))  severity failure;
	assert RAM(18551) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(18551))))  severity failure;
	assert RAM(18552) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(18552))))  severity failure;
	assert RAM(18553) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(18553))))  severity failure;
	assert RAM(18554) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(18554))))  severity failure;
	assert RAM(18555) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(18555))))  severity failure;
	assert RAM(18556) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(18556))))  severity failure;
	assert RAM(18557) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(18557))))  severity failure;
	assert RAM(18558) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(18558))))  severity failure;
	assert RAM(18559) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(18559))))  severity failure;
	assert RAM(18560) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(18560))))  severity failure;
	assert RAM(18561) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18561))))  severity failure;
	assert RAM(18562) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18562))))  severity failure;
	assert RAM(18563) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(18563))))  severity failure;
	assert RAM(18564) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18564))))  severity failure;
	assert RAM(18565) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(18565))))  severity failure;
	assert RAM(18566) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(18566))))  severity failure;
	assert RAM(18567) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(18567))))  severity failure;
	assert RAM(18568) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18568))))  severity failure;
	assert RAM(18569) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(18569))))  severity failure;
	assert RAM(18570) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(18570))))  severity failure;
	assert RAM(18571) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(18571))))  severity failure;
	assert RAM(18572) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(18572))))  severity failure;
	assert RAM(18573) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18573))))  severity failure;
	assert RAM(18574) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(18574))))  severity failure;
	assert RAM(18575) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18575))))  severity failure;
	assert RAM(18576) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(18576))))  severity failure;
	assert RAM(18577) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(18577))))  severity failure;
	assert RAM(18578) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(18578))))  severity failure;
	assert RAM(18579) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(18579))))  severity failure;
	assert RAM(18580) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(18580))))  severity failure;
	assert RAM(18581) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(18581))))  severity failure;
	assert RAM(18582) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(18582))))  severity failure;
	assert RAM(18583) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(18583))))  severity failure;
	assert RAM(18584) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(18584))))  severity failure;
	assert RAM(18585) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18585))))  severity failure;
	assert RAM(18586) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(18586))))  severity failure;
	assert RAM(18587) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(18587))))  severity failure;
	assert RAM(18588) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(18588))))  severity failure;
	assert RAM(18589) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(18589))))  severity failure;
	assert RAM(18590) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18590))))  severity failure;
	assert RAM(18591) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(18591))))  severity failure;
	assert RAM(18592) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(18592))))  severity failure;
	assert RAM(18593) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(18593))))  severity failure;
	assert RAM(18594) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(18594))))  severity failure;
	assert RAM(18595) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(18595))))  severity failure;
	assert RAM(18596) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18596))))  severity failure;
	assert RAM(18597) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(18597))))  severity failure;
	assert RAM(18598) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18598))))  severity failure;
	assert RAM(18599) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18599))))  severity failure;
	assert RAM(18600) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(18600))))  severity failure;
	assert RAM(18601) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(18601))))  severity failure;
	assert RAM(18602) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(18602))))  severity failure;
	assert RAM(18603) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18603))))  severity failure;
	assert RAM(18604) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(18604))))  severity failure;
	assert RAM(18605) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(18605))))  severity failure;
	assert RAM(18606) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(18606))))  severity failure;
	assert RAM(18607) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18607))))  severity failure;
	assert RAM(18608) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(18608))))  severity failure;
	assert RAM(18609) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18609))))  severity failure;
	assert RAM(18610) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(18610))))  severity failure;
	assert RAM(18611) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18611))))  severity failure;
	assert RAM(18612) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(18612))))  severity failure;
	assert RAM(18613) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(18613))))  severity failure;
	assert RAM(18614) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(18614))))  severity failure;
	assert RAM(18615) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18615))))  severity failure;
	assert RAM(18616) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18616))))  severity failure;
	assert RAM(18617) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(18617))))  severity failure;
	assert RAM(18618) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(18618))))  severity failure;
	assert RAM(18619) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(18619))))  severity failure;
	assert RAM(18620) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(18620))))  severity failure;
	assert RAM(18621) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(18621))))  severity failure;
	assert RAM(18622) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(18622))))  severity failure;
	assert RAM(18623) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(18623))))  severity failure;
	assert RAM(18624) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(18624))))  severity failure;
	assert RAM(18625) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(18625))))  severity failure;
	assert RAM(18626) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(18626))))  severity failure;
	assert RAM(18627) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18627))))  severity failure;
	assert RAM(18628) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18628))))  severity failure;
	assert RAM(18629) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18629))))  severity failure;
	assert RAM(18630) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(18630))))  severity failure;
	assert RAM(18631) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(18631))))  severity failure;
	assert RAM(18632) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(18632))))  severity failure;
	assert RAM(18633) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(18633))))  severity failure;
	assert RAM(18634) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(18634))))  severity failure;
	assert RAM(18635) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18635))))  severity failure;
	assert RAM(18636) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(18636))))  severity failure;
	assert RAM(18637) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(18637))))  severity failure;
	assert RAM(18638) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18638))))  severity failure;
	assert RAM(18639) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(18639))))  severity failure;
	assert RAM(18640) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(18640))))  severity failure;
	assert RAM(18641) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(18641))))  severity failure;
	assert RAM(18642) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(18642))))  severity failure;
	assert RAM(18643) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(18643))))  severity failure;
	assert RAM(18644) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(18644))))  severity failure;
	assert RAM(18645) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18645))))  severity failure;
	assert RAM(18646) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(18646))))  severity failure;
	assert RAM(18647) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(18647))))  severity failure;
	assert RAM(18648) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18648))))  severity failure;
	assert RAM(18649) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(18649))))  severity failure;
	assert RAM(18650) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(18650))))  severity failure;
	assert RAM(18651) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(18651))))  severity failure;
	assert RAM(18652) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(18652))))  severity failure;
	assert RAM(18653) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18653))))  severity failure;
	assert RAM(18654) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18654))))  severity failure;
	assert RAM(18655) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(18655))))  severity failure;
	assert RAM(18656) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(18656))))  severity failure;
	assert RAM(18657) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(18657))))  severity failure;
	assert RAM(18658) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(18658))))  severity failure;
	assert RAM(18659) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(18659))))  severity failure;
	assert RAM(18660) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18660))))  severity failure;
	assert RAM(18661) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(18661))))  severity failure;
	assert RAM(18662) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(18662))))  severity failure;
	assert RAM(18663) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(18663))))  severity failure;
	assert RAM(18664) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18664))))  severity failure;
	assert RAM(18665) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18665))))  severity failure;
	assert RAM(18666) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(18666))))  severity failure;
	assert RAM(18667) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(18667))))  severity failure;
	assert RAM(18668) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(18668))))  severity failure;
	assert RAM(18669) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(18669))))  severity failure;
	assert RAM(18670) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(18670))))  severity failure;
	assert RAM(18671) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18671))))  severity failure;
	assert RAM(18672) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(18672))))  severity failure;
	assert RAM(18673) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(18673))))  severity failure;
	assert RAM(18674) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(18674))))  severity failure;
	assert RAM(18675) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(18675))))  severity failure;
	assert RAM(18676) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(18676))))  severity failure;
	assert RAM(18677) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(18677))))  severity failure;
	assert RAM(18678) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(18678))))  severity failure;
	assert RAM(18679) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(18679))))  severity failure;
	assert RAM(18680) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(18680))))  severity failure;
	assert RAM(18681) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(18681))))  severity failure;
	assert RAM(18682) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(18682))))  severity failure;
	assert RAM(18683) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(18683))))  severity failure;
	assert RAM(18684) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(18684))))  severity failure;
	assert RAM(18685) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(18685))))  severity failure;
	assert RAM(18686) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(18686))))  severity failure;
	assert RAM(18687) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(18687))))  severity failure;
	assert RAM(18688) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18688))))  severity failure;
	assert RAM(18689) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(18689))))  severity failure;
	assert RAM(18690) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(18690))))  severity failure;
	assert RAM(18691) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(18691))))  severity failure;
	assert RAM(18692) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(18692))))  severity failure;
	assert RAM(18693) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(18693))))  severity failure;
	assert RAM(18694) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(18694))))  severity failure;
	assert RAM(18695) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(18695))))  severity failure;
	assert RAM(18696) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(18696))))  severity failure;
	assert RAM(18697) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(18697))))  severity failure;
	assert RAM(18698) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(18698))))  severity failure;
	assert RAM(18699) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(18699))))  severity failure;
	assert RAM(18700) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(18700))))  severity failure;
	assert RAM(18701) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(18701))))  severity failure;
	assert RAM(18702) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(18702))))  severity failure;
	assert RAM(18703) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(18703))))  severity failure;
	assert RAM(18704) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(18704))))  severity failure;
	assert RAM(18705) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18705))))  severity failure;
	assert RAM(18706) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(18706))))  severity failure;
	assert RAM(18707) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(18707))))  severity failure;
	assert RAM(18708) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(18708))))  severity failure;
	assert RAM(18709) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(18709))))  severity failure;
	assert RAM(18710) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(18710))))  severity failure;
	assert RAM(18711) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(18711))))  severity failure;
	assert RAM(18712) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(18712))))  severity failure;
	assert RAM(18713) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18713))))  severity failure;
	assert RAM(18714) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(18714))))  severity failure;
	assert RAM(18715) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(18715))))  severity failure;
	assert RAM(18716) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18716))))  severity failure;
	assert RAM(18717) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(18717))))  severity failure;
	assert RAM(18718) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18718))))  severity failure;
	assert RAM(18719) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(18719))))  severity failure;
	assert RAM(18720) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(18720))))  severity failure;
	assert RAM(18721) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(18721))))  severity failure;
	assert RAM(18722) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(18722))))  severity failure;
	assert RAM(18723) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(18723))))  severity failure;
	assert RAM(18724) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18724))))  severity failure;
	assert RAM(18725) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18725))))  severity failure;
	assert RAM(18726) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(18726))))  severity failure;
	assert RAM(18727) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18727))))  severity failure;
	assert RAM(18728) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(18728))))  severity failure;
	assert RAM(18729) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(18729))))  severity failure;
	assert RAM(18730) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(18730))))  severity failure;
	assert RAM(18731) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(18731))))  severity failure;
	assert RAM(18732) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(18732))))  severity failure;
	assert RAM(18733) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(18733))))  severity failure;
	assert RAM(18734) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18734))))  severity failure;
	assert RAM(18735) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18735))))  severity failure;
	assert RAM(18736) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(18736))))  severity failure;
	assert RAM(18737) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(18737))))  severity failure;
	assert RAM(18738) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(18738))))  severity failure;
	assert RAM(18739) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(18739))))  severity failure;
	assert RAM(18740) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18740))))  severity failure;
	assert RAM(18741) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(18741))))  severity failure;
	assert RAM(18742) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(18742))))  severity failure;
	assert RAM(18743) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18743))))  severity failure;
	assert RAM(18744) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18744))))  severity failure;
	assert RAM(18745) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(18745))))  severity failure;
	assert RAM(18746) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(18746))))  severity failure;
	assert RAM(18747) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18747))))  severity failure;
	assert RAM(18748) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(18748))))  severity failure;
	assert RAM(18749) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18749))))  severity failure;
	assert RAM(18750) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(18750))))  severity failure;
	assert RAM(18751) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(18751))))  severity failure;
	assert RAM(18752) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(18752))))  severity failure;
	assert RAM(18753) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(18753))))  severity failure;
	assert RAM(18754) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(18754))))  severity failure;
	assert RAM(18755) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(18755))))  severity failure;
	assert RAM(18756) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(18756))))  severity failure;
	assert RAM(18757) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18757))))  severity failure;
	assert RAM(18758) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(18758))))  severity failure;
	assert RAM(18759) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(18759))))  severity failure;
	assert RAM(18760) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18760))))  severity failure;
	assert RAM(18761) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(18761))))  severity failure;
	assert RAM(18762) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18762))))  severity failure;
	assert RAM(18763) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(18763))))  severity failure;
	assert RAM(18764) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(18764))))  severity failure;
	assert RAM(18765) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(18765))))  severity failure;
	assert RAM(18766) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18766))))  severity failure;
	assert RAM(18767) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(18767))))  severity failure;
	assert RAM(18768) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18768))))  severity failure;
	assert RAM(18769) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(18769))))  severity failure;
	assert RAM(18770) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18770))))  severity failure;
	assert RAM(18771) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(18771))))  severity failure;
	assert RAM(18772) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(18772))))  severity failure;
	assert RAM(18773) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(18773))))  severity failure;
	assert RAM(18774) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(18774))))  severity failure;
	assert RAM(18775) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(18775))))  severity failure;
	assert RAM(18776) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18776))))  severity failure;
	assert RAM(18777) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(18777))))  severity failure;
	assert RAM(18778) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(18778))))  severity failure;
	assert RAM(18779) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(18779))))  severity failure;
	assert RAM(18780) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18780))))  severity failure;
	assert RAM(18781) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(18781))))  severity failure;
	assert RAM(18782) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18782))))  severity failure;
	assert RAM(18783) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(18783))))  severity failure;
	assert RAM(18784) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(18784))))  severity failure;
	assert RAM(18785) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(18785))))  severity failure;
	assert RAM(18786) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18786))))  severity failure;
	assert RAM(18787) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(18787))))  severity failure;
	assert RAM(18788) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(18788))))  severity failure;
	assert RAM(18789) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18789))))  severity failure;
	assert RAM(18790) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18790))))  severity failure;
	assert RAM(18791) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18791))))  severity failure;
	assert RAM(18792) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18792))))  severity failure;
	assert RAM(18793) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(18793))))  severity failure;
	assert RAM(18794) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(18794))))  severity failure;
	assert RAM(18795) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(18795))))  severity failure;
	assert RAM(18796) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(18796))))  severity failure;
	assert RAM(18797) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(18797))))  severity failure;
	assert RAM(18798) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18798))))  severity failure;
	assert RAM(18799) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(18799))))  severity failure;
	assert RAM(18800) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18800))))  severity failure;
	assert RAM(18801) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(18801))))  severity failure;
	assert RAM(18802) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(18802))))  severity failure;
	assert RAM(18803) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18803))))  severity failure;
	assert RAM(18804) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(18804))))  severity failure;
	assert RAM(18805) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(18805))))  severity failure;
	assert RAM(18806) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(18806))))  severity failure;
	assert RAM(18807) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18807))))  severity failure;
	assert RAM(18808) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(18808))))  severity failure;
	assert RAM(18809) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(18809))))  severity failure;
	assert RAM(18810) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(18810))))  severity failure;
	assert RAM(18811) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18811))))  severity failure;
	assert RAM(18812) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18812))))  severity failure;
	assert RAM(18813) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(18813))))  severity failure;
	assert RAM(18814) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(18814))))  severity failure;
	assert RAM(18815) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(18815))))  severity failure;
	assert RAM(18816) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(18816))))  severity failure;
	assert RAM(18817) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(18817))))  severity failure;
	assert RAM(18818) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18818))))  severity failure;
	assert RAM(18819) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(18819))))  severity failure;
	assert RAM(18820) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18820))))  severity failure;
	assert RAM(18821) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(18821))))  severity failure;
	assert RAM(18822) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(18822))))  severity failure;
	assert RAM(18823) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(18823))))  severity failure;
	assert RAM(18824) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(18824))))  severity failure;
	assert RAM(18825) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(18825))))  severity failure;
	assert RAM(18826) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(18826))))  severity failure;
	assert RAM(18827) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18827))))  severity failure;
	assert RAM(18828) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(18828))))  severity failure;
	assert RAM(18829) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(18829))))  severity failure;
	assert RAM(18830) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18830))))  severity failure;
	assert RAM(18831) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18831))))  severity failure;
	assert RAM(18832) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(18832))))  severity failure;
	assert RAM(18833) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(18833))))  severity failure;
	assert RAM(18834) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18834))))  severity failure;
	assert RAM(18835) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18835))))  severity failure;
	assert RAM(18836) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(18836))))  severity failure;
	assert RAM(18837) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(18837))))  severity failure;
	assert RAM(18838) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(18838))))  severity failure;
	assert RAM(18839) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(18839))))  severity failure;
	assert RAM(18840) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(18840))))  severity failure;
	assert RAM(18841) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18841))))  severity failure;
	assert RAM(18842) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(18842))))  severity failure;
	assert RAM(18843) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(18843))))  severity failure;
	assert RAM(18844) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(18844))))  severity failure;
	assert RAM(18845) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18845))))  severity failure;
	assert RAM(18846) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(18846))))  severity failure;
	assert RAM(18847) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(18847))))  severity failure;
	assert RAM(18848) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(18848))))  severity failure;
	assert RAM(18849) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(18849))))  severity failure;
	assert RAM(18850) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(18850))))  severity failure;
	assert RAM(18851) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(18851))))  severity failure;
	assert RAM(18852) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(18852))))  severity failure;
	assert RAM(18853) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(18853))))  severity failure;
	assert RAM(18854) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(18854))))  severity failure;
	assert RAM(18855) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(18855))))  severity failure;
	assert RAM(18856) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(18856))))  severity failure;
	assert RAM(18857) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(18857))))  severity failure;
	assert RAM(18858) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(18858))))  severity failure;
	assert RAM(18859) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(18859))))  severity failure;
	assert RAM(18860) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(18860))))  severity failure;
	assert RAM(18861) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18861))))  severity failure;
	assert RAM(18862) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(18862))))  severity failure;
	assert RAM(18863) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(18863))))  severity failure;
	assert RAM(18864) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(18864))))  severity failure;
	assert RAM(18865) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18865))))  severity failure;
	assert RAM(18866) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(18866))))  severity failure;
	assert RAM(18867) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(18867))))  severity failure;
	assert RAM(18868) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18868))))  severity failure;
	assert RAM(18869) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(18869))))  severity failure;
	assert RAM(18870) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(18870))))  severity failure;
	assert RAM(18871) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(18871))))  severity failure;
	assert RAM(18872) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18872))))  severity failure;
	assert RAM(18873) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18873))))  severity failure;
	assert RAM(18874) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(18874))))  severity failure;
	assert RAM(18875) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(18875))))  severity failure;
	assert RAM(18876) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(18876))))  severity failure;
	assert RAM(18877) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(18877))))  severity failure;
	assert RAM(18878) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(18878))))  severity failure;
	assert RAM(18879) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(18879))))  severity failure;
	assert RAM(18880) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(18880))))  severity failure;
	assert RAM(18881) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(18881))))  severity failure;
	assert RAM(18882) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18882))))  severity failure;
	assert RAM(18883) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(18883))))  severity failure;
	assert RAM(18884) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(18884))))  severity failure;
	assert RAM(18885) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(18885))))  severity failure;
	assert RAM(18886) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(18886))))  severity failure;
	assert RAM(18887) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(18887))))  severity failure;
	assert RAM(18888) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18888))))  severity failure;
	assert RAM(18889) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(18889))))  severity failure;
	assert RAM(18890) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(18890))))  severity failure;
	assert RAM(18891) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(18891))))  severity failure;
	assert RAM(18892) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(18892))))  severity failure;
	assert RAM(18893) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(18893))))  severity failure;
	assert RAM(18894) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(18894))))  severity failure;
	assert RAM(18895) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(18895))))  severity failure;
	assert RAM(18896) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(18896))))  severity failure;
	assert RAM(18897) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(18897))))  severity failure;
	assert RAM(18898) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18898))))  severity failure;
	assert RAM(18899) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(18899))))  severity failure;
	assert RAM(18900) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(18900))))  severity failure;
	assert RAM(18901) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18901))))  severity failure;
	assert RAM(18902) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(18902))))  severity failure;
	assert RAM(18903) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(18903))))  severity failure;
	assert RAM(18904) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(18904))))  severity failure;
	assert RAM(18905) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(18905))))  severity failure;
	assert RAM(18906) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(18906))))  severity failure;
	assert RAM(18907) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(18907))))  severity failure;
	assert RAM(18908) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(18908))))  severity failure;
	assert RAM(18909) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(18909))))  severity failure;
	assert RAM(18910) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(18910))))  severity failure;
	assert RAM(18911) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18911))))  severity failure;
	assert RAM(18912) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(18912))))  severity failure;
	assert RAM(18913) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(18913))))  severity failure;
	assert RAM(18914) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(18914))))  severity failure;
	assert RAM(18915) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(18915))))  severity failure;
	assert RAM(18916) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18916))))  severity failure;
	assert RAM(18917) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18917))))  severity failure;
	assert RAM(18918) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(18918))))  severity failure;
	assert RAM(18919) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(18919))))  severity failure;
	assert RAM(18920) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(18920))))  severity failure;
	assert RAM(18921) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(18921))))  severity failure;
	assert RAM(18922) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(18922))))  severity failure;
	assert RAM(18923) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(18923))))  severity failure;
	assert RAM(18924) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18924))))  severity failure;
	assert RAM(18925) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(18925))))  severity failure;
	assert RAM(18926) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(18926))))  severity failure;
	assert RAM(18927) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(18927))))  severity failure;
	assert RAM(18928) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(18928))))  severity failure;
	assert RAM(18929) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18929))))  severity failure;
	assert RAM(18930) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(18930))))  severity failure;
	assert RAM(18931) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18931))))  severity failure;
	assert RAM(18932) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(18932))))  severity failure;
	assert RAM(18933) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(18933))))  severity failure;
	assert RAM(18934) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(18934))))  severity failure;
	assert RAM(18935) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18935))))  severity failure;
	assert RAM(18936) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(18936))))  severity failure;
	assert RAM(18937) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(18937))))  severity failure;
	assert RAM(18938) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(18938))))  severity failure;
	assert RAM(18939) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(18939))))  severity failure;
	assert RAM(18940) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(18940))))  severity failure;
	assert RAM(18941) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(18941))))  severity failure;
	assert RAM(18942) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(18942))))  severity failure;
	assert RAM(18943) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(18943))))  severity failure;
	assert RAM(18944) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(18944))))  severity failure;
	assert RAM(18945) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(18945))))  severity failure;
	assert RAM(18946) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(18946))))  severity failure;
	assert RAM(18947) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(18947))))  severity failure;
	assert RAM(18948) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(18948))))  severity failure;
	assert RAM(18949) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(18949))))  severity failure;
	assert RAM(18950) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(18950))))  severity failure;
	assert RAM(18951) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(18951))))  severity failure;
	assert RAM(18952) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(18952))))  severity failure;
	assert RAM(18953) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(18953))))  severity failure;
	assert RAM(18954) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(18954))))  severity failure;
	assert RAM(18955) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(18955))))  severity failure;
	assert RAM(18956) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(18956))))  severity failure;
	assert RAM(18957) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(18957))))  severity failure;
	assert RAM(18958) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(18958))))  severity failure;
	assert RAM(18959) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(18959))))  severity failure;
	assert RAM(18960) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(18960))))  severity failure;
	assert RAM(18961) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(18961))))  severity failure;
	assert RAM(18962) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(18962))))  severity failure;
	assert RAM(18963) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(18963))))  severity failure;
	assert RAM(18964) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(18964))))  severity failure;
	assert RAM(18965) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(18965))))  severity failure;
	assert RAM(18966) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(18966))))  severity failure;
	assert RAM(18967) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(18967))))  severity failure;
	assert RAM(18968) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(18968))))  severity failure;
	assert RAM(18969) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(18969))))  severity failure;
	assert RAM(18970) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(18970))))  severity failure;
	assert RAM(18971) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(18971))))  severity failure;
	assert RAM(18972) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(18972))))  severity failure;
	assert RAM(18973) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(18973))))  severity failure;
	assert RAM(18974) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(18974))))  severity failure;
	assert RAM(18975) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(18975))))  severity failure;
	assert RAM(18976) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(18976))))  severity failure;
	assert RAM(18977) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(18977))))  severity failure;
	assert RAM(18978) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(18978))))  severity failure;
	assert RAM(18979) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(18979))))  severity failure;
	assert RAM(18980) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(18980))))  severity failure;
	assert RAM(18981) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(18981))))  severity failure;
	assert RAM(18982) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(18982))))  severity failure;
	assert RAM(18983) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(18983))))  severity failure;
	assert RAM(18984) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(18984))))  severity failure;
	assert RAM(18985) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(18985))))  severity failure;
	assert RAM(18986) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(18986))))  severity failure;
	assert RAM(18987) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(18987))))  severity failure;
	assert RAM(18988) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(18988))))  severity failure;
	assert RAM(18989) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(18989))))  severity failure;
	assert RAM(18990) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(18990))))  severity failure;
	assert RAM(18991) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(18991))))  severity failure;
	assert RAM(18992) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(18992))))  severity failure;
	assert RAM(18993) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(18993))))  severity failure;
	assert RAM(18994) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(18994))))  severity failure;
	assert RAM(18995) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(18995))))  severity failure;
	assert RAM(18996) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(18996))))  severity failure;
	assert RAM(18997) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(18997))))  severity failure;
	assert RAM(18998) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(18998))))  severity failure;
	assert RAM(18999) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(18999))))  severity failure;
	assert RAM(19000) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19000))))  severity failure;
	assert RAM(19001) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(19001))))  severity failure;
	assert RAM(19002) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19002))))  severity failure;
	assert RAM(19003) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(19003))))  severity failure;
	assert RAM(19004) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(19004))))  severity failure;
	assert RAM(19005) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19005))))  severity failure;
	assert RAM(19006) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19006))))  severity failure;
	assert RAM(19007) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19007))))  severity failure;
	assert RAM(19008) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19008))))  severity failure;
	assert RAM(19009) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(19009))))  severity failure;
	assert RAM(19010) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(19010))))  severity failure;
	assert RAM(19011) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19011))))  severity failure;
	assert RAM(19012) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(19012))))  severity failure;
	assert RAM(19013) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(19013))))  severity failure;
	assert RAM(19014) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(19014))))  severity failure;
	assert RAM(19015) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19015))))  severity failure;
	assert RAM(19016) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(19016))))  severity failure;
	assert RAM(19017) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(19017))))  severity failure;
	assert RAM(19018) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19018))))  severity failure;
	assert RAM(19019) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19019))))  severity failure;
	assert RAM(19020) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19020))))  severity failure;
	assert RAM(19021) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(19021))))  severity failure;
	assert RAM(19022) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(19022))))  severity failure;
	assert RAM(19023) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(19023))))  severity failure;
	assert RAM(19024) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(19024))))  severity failure;
	assert RAM(19025) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(19025))))  severity failure;
	assert RAM(19026) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(19026))))  severity failure;
	assert RAM(19027) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(19027))))  severity failure;
	assert RAM(19028) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(19028))))  severity failure;
	assert RAM(19029) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(19029))))  severity failure;
	assert RAM(19030) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(19030))))  severity failure;
	assert RAM(19031) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(19031))))  severity failure;
	assert RAM(19032) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(19032))))  severity failure;
	assert RAM(19033) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19033))))  severity failure;
	assert RAM(19034) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(19034))))  severity failure;
	assert RAM(19035) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(19035))))  severity failure;
	assert RAM(19036) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(19036))))  severity failure;
	assert RAM(19037) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19037))))  severity failure;
	assert RAM(19038) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(19038))))  severity failure;
	assert RAM(19039) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(19039))))  severity failure;
	assert RAM(19040) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19040))))  severity failure;
	assert RAM(19041) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(19041))))  severity failure;
	assert RAM(19042) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(19042))))  severity failure;
	assert RAM(19043) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19043))))  severity failure;
	assert RAM(19044) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(19044))))  severity failure;
	assert RAM(19045) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(19045))))  severity failure;
	assert RAM(19046) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(19046))))  severity failure;
	assert RAM(19047) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(19047))))  severity failure;
	assert RAM(19048) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19048))))  severity failure;
	assert RAM(19049) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(19049))))  severity failure;
	assert RAM(19050) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(19050))))  severity failure;
	assert RAM(19051) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19051))))  severity failure;
	assert RAM(19052) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19052))))  severity failure;
	assert RAM(19053) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(19053))))  severity failure;
	assert RAM(19054) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(19054))))  severity failure;
	assert RAM(19055) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(19055))))  severity failure;
	assert RAM(19056) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(19056))))  severity failure;
	assert RAM(19057) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19057))))  severity failure;
	assert RAM(19058) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(19058))))  severity failure;
	assert RAM(19059) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(19059))))  severity failure;
	assert RAM(19060) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(19060))))  severity failure;
	assert RAM(19061) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19061))))  severity failure;
	assert RAM(19062) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(19062))))  severity failure;
	assert RAM(19063) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(19063))))  severity failure;
	assert RAM(19064) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(19064))))  severity failure;
	assert RAM(19065) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(19065))))  severity failure;
	assert RAM(19066) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(19066))))  severity failure;
	assert RAM(19067) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(19067))))  severity failure;
	assert RAM(19068) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(19068))))  severity failure;
	assert RAM(19069) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(19069))))  severity failure;
	assert RAM(19070) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19070))))  severity failure;
	assert RAM(19071) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(19071))))  severity failure;
	assert RAM(19072) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(19072))))  severity failure;
	assert RAM(19073) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(19073))))  severity failure;
	assert RAM(19074) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(19074))))  severity failure;
	assert RAM(19075) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(19075))))  severity failure;
	assert RAM(19076) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(19076))))  severity failure;
	assert RAM(19077) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(19077))))  severity failure;
	assert RAM(19078) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(19078))))  severity failure;
	assert RAM(19079) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(19079))))  severity failure;
	assert RAM(19080) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(19080))))  severity failure;
	assert RAM(19081) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19081))))  severity failure;
	assert RAM(19082) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(19082))))  severity failure;
	assert RAM(19083) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(19083))))  severity failure;
	assert RAM(19084) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(19084))))  severity failure;
	assert RAM(19085) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(19085))))  severity failure;
	assert RAM(19086) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(19086))))  severity failure;
	assert RAM(19087) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19087))))  severity failure;
	assert RAM(19088) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(19088))))  severity failure;
	assert RAM(19089) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(19089))))  severity failure;
	assert RAM(19090) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(19090))))  severity failure;
	assert RAM(19091) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(19091))))  severity failure;
	assert RAM(19092) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19092))))  severity failure;
	assert RAM(19093) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19093))))  severity failure;
	assert RAM(19094) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(19094))))  severity failure;
	assert RAM(19095) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(19095))))  severity failure;
	assert RAM(19096) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19096))))  severity failure;
	assert RAM(19097) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19097))))  severity failure;
	assert RAM(19098) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(19098))))  severity failure;
	assert RAM(19099) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(19099))))  severity failure;
	assert RAM(19100) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19100))))  severity failure;
	assert RAM(19101) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19101))))  severity failure;
	assert RAM(19102) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(19102))))  severity failure;
	assert RAM(19103) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(19103))))  severity failure;
	assert RAM(19104) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19104))))  severity failure;
	assert RAM(19105) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(19105))))  severity failure;
	assert RAM(19106) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(19106))))  severity failure;
	assert RAM(19107) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19107))))  severity failure;
	assert RAM(19108) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(19108))))  severity failure;
	assert RAM(19109) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(19109))))  severity failure;
	assert RAM(19110) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(19110))))  severity failure;
	assert RAM(19111) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(19111))))  severity failure;
	assert RAM(19112) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(19112))))  severity failure;
	assert RAM(19113) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19113))))  severity failure;
	assert RAM(19114) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(19114))))  severity failure;
	assert RAM(19115) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(19115))))  severity failure;
	assert RAM(19116) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(19116))))  severity failure;
	assert RAM(19117) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19117))))  severity failure;
	assert RAM(19118) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19118))))  severity failure;
	assert RAM(19119) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(19119))))  severity failure;
	assert RAM(19120) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19120))))  severity failure;
	assert RAM(19121) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(19121))))  severity failure;
	assert RAM(19122) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(19122))))  severity failure;
	assert RAM(19123) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(19123))))  severity failure;
	assert RAM(19124) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(19124))))  severity failure;
	assert RAM(19125) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(19125))))  severity failure;
	assert RAM(19126) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(19126))))  severity failure;
	assert RAM(19127) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(19127))))  severity failure;
	assert RAM(19128) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(19128))))  severity failure;
	assert RAM(19129) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19129))))  severity failure;
	assert RAM(19130) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19130))))  severity failure;
	assert RAM(19131) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(19131))))  severity failure;
	assert RAM(19132) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(19132))))  severity failure;
	assert RAM(19133) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19133))))  severity failure;
	assert RAM(19134) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(19134))))  severity failure;
	assert RAM(19135) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(19135))))  severity failure;
	assert RAM(19136) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19136))))  severity failure;
	assert RAM(19137) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(19137))))  severity failure;
	assert RAM(19138) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19138))))  severity failure;
	assert RAM(19139) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19139))))  severity failure;
	assert RAM(19140) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19140))))  severity failure;
	assert RAM(19141) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19141))))  severity failure;
	assert RAM(19142) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(19142))))  severity failure;
	assert RAM(19143) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(19143))))  severity failure;
	assert RAM(19144) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19144))))  severity failure;
	assert RAM(19145) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(19145))))  severity failure;
	assert RAM(19146) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(19146))))  severity failure;
	assert RAM(19147) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19147))))  severity failure;
	assert RAM(19148) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(19148))))  severity failure;
	assert RAM(19149) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(19149))))  severity failure;
	assert RAM(19150) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19150))))  severity failure;
	assert RAM(19151) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(19151))))  severity failure;
	assert RAM(19152) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(19152))))  severity failure;
	assert RAM(19153) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(19153))))  severity failure;
	assert RAM(19154) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(19154))))  severity failure;
	assert RAM(19155) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(19155))))  severity failure;
	assert RAM(19156) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19156))))  severity failure;
	assert RAM(19157) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19157))))  severity failure;
	assert RAM(19158) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(19158))))  severity failure;
	assert RAM(19159) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(19159))))  severity failure;
	assert RAM(19160) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(19160))))  severity failure;
	assert RAM(19161) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19161))))  severity failure;
	assert RAM(19162) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(19162))))  severity failure;
	assert RAM(19163) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(19163))))  severity failure;
	assert RAM(19164) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(19164))))  severity failure;
	assert RAM(19165) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(19165))))  severity failure;
	assert RAM(19166) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19166))))  severity failure;
	assert RAM(19167) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(19167))))  severity failure;
	assert RAM(19168) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(19168))))  severity failure;
	assert RAM(19169) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19169))))  severity failure;
	assert RAM(19170) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(19170))))  severity failure;
	assert RAM(19171) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19171))))  severity failure;
	assert RAM(19172) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19172))))  severity failure;
	assert RAM(19173) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(19173))))  severity failure;
	assert RAM(19174) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(19174))))  severity failure;
	assert RAM(19175) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(19175))))  severity failure;
	assert RAM(19176) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(19176))))  severity failure;
	assert RAM(19177) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(19177))))  severity failure;
	assert RAM(19178) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19178))))  severity failure;
	assert RAM(19179) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(19179))))  severity failure;
	assert RAM(19180) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(19180))))  severity failure;
	assert RAM(19181) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(19181))))  severity failure;
	assert RAM(19182) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(19182))))  severity failure;
	assert RAM(19183) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(19183))))  severity failure;
	assert RAM(19184) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(19184))))  severity failure;
	assert RAM(19185) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(19185))))  severity failure;
	assert RAM(19186) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(19186))))  severity failure;
	assert RAM(19187) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19187))))  severity failure;
	assert RAM(19188) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(19188))))  severity failure;
	assert RAM(19189) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(19189))))  severity failure;
	assert RAM(19190) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(19190))))  severity failure;
	assert RAM(19191) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(19191))))  severity failure;
	assert RAM(19192) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(19192))))  severity failure;
	assert RAM(19193) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(19193))))  severity failure;
	assert RAM(19194) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(19194))))  severity failure;
	assert RAM(19195) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19195))))  severity failure;
	assert RAM(19196) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19196))))  severity failure;
	assert RAM(19197) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(19197))))  severity failure;
	assert RAM(19198) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(19198))))  severity failure;
	assert RAM(19199) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19199))))  severity failure;
	assert RAM(19200) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(19200))))  severity failure;
	assert RAM(19201) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(19201))))  severity failure;
	assert RAM(19202) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(19202))))  severity failure;
	assert RAM(19203) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(19203))))  severity failure;
	assert RAM(19204) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(19204))))  severity failure;
	assert RAM(19205) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19205))))  severity failure;
	assert RAM(19206) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(19206))))  severity failure;
	assert RAM(19207) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19207))))  severity failure;
	assert RAM(19208) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(19208))))  severity failure;
	assert RAM(19209) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19209))))  severity failure;
	assert RAM(19210) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19210))))  severity failure;
	assert RAM(19211) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19211))))  severity failure;
	assert RAM(19212) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(19212))))  severity failure;
	assert RAM(19213) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(19213))))  severity failure;
	assert RAM(19214) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(19214))))  severity failure;
	assert RAM(19215) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(19215))))  severity failure;
	assert RAM(19216) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(19216))))  severity failure;
	assert RAM(19217) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(19217))))  severity failure;
	assert RAM(19218) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(19218))))  severity failure;
	assert RAM(19219) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(19219))))  severity failure;
	assert RAM(19220) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(19220))))  severity failure;
	assert RAM(19221) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(19221))))  severity failure;
	assert RAM(19222) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(19222))))  severity failure;
	assert RAM(19223) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19223))))  severity failure;
	assert RAM(19224) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(19224))))  severity failure;
	assert RAM(19225) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19225))))  severity failure;
	assert RAM(19226) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(19226))))  severity failure;
	assert RAM(19227) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19227))))  severity failure;
	assert RAM(19228) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19228))))  severity failure;
	assert RAM(19229) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(19229))))  severity failure;
	assert RAM(19230) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(19230))))  severity failure;
	assert RAM(19231) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(19231))))  severity failure;
	assert RAM(19232) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19232))))  severity failure;
	assert RAM(19233) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(19233))))  severity failure;
	assert RAM(19234) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(19234))))  severity failure;
	assert RAM(19235) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19235))))  severity failure;
	assert RAM(19236) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(19236))))  severity failure;
	assert RAM(19237) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19237))))  severity failure;
	assert RAM(19238) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(19238))))  severity failure;
	assert RAM(19239) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19239))))  severity failure;
	assert RAM(19240) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(19240))))  severity failure;
	assert RAM(19241) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(19241))))  severity failure;
	assert RAM(19242) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(19242))))  severity failure;
	assert RAM(19243) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(19243))))  severity failure;
	assert RAM(19244) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(19244))))  severity failure;
	assert RAM(19245) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(19245))))  severity failure;
	assert RAM(19246) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(19246))))  severity failure;
	assert RAM(19247) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19247))))  severity failure;
	assert RAM(19248) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(19248))))  severity failure;
	assert RAM(19249) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(19249))))  severity failure;
	assert RAM(19250) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(19250))))  severity failure;
	assert RAM(19251) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19251))))  severity failure;
	assert RAM(19252) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(19252))))  severity failure;
	assert RAM(19253) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(19253))))  severity failure;
	assert RAM(19254) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(19254))))  severity failure;
	assert RAM(19255) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(19255))))  severity failure;
	assert RAM(19256) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(19256))))  severity failure;
	assert RAM(19257) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(19257))))  severity failure;
	assert RAM(19258) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(19258))))  severity failure;
	assert RAM(19259) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(19259))))  severity failure;
	assert RAM(19260) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19260))))  severity failure;
	assert RAM(19261) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19261))))  severity failure;
	assert RAM(19262) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(19262))))  severity failure;
	assert RAM(19263) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(19263))))  severity failure;
	assert RAM(19264) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19264))))  severity failure;
	assert RAM(19265) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(19265))))  severity failure;
	assert RAM(19266) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(19266))))  severity failure;
	assert RAM(19267) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(19267))))  severity failure;
	assert RAM(19268) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19268))))  severity failure;
	assert RAM(19269) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(19269))))  severity failure;
	assert RAM(19270) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(19270))))  severity failure;
	assert RAM(19271) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19271))))  severity failure;
	assert RAM(19272) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(19272))))  severity failure;
	assert RAM(19273) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(19273))))  severity failure;
	assert RAM(19274) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(19274))))  severity failure;
	assert RAM(19275) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(19275))))  severity failure;
	assert RAM(19276) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(19276))))  severity failure;
	assert RAM(19277) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19277))))  severity failure;
	assert RAM(19278) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19278))))  severity failure;
	assert RAM(19279) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(19279))))  severity failure;
	assert RAM(19280) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(19280))))  severity failure;
	assert RAM(19281) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(19281))))  severity failure;
	assert RAM(19282) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(19282))))  severity failure;
	assert RAM(19283) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(19283))))  severity failure;
	assert RAM(19284) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(19284))))  severity failure;
	assert RAM(19285) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19285))))  severity failure;
	assert RAM(19286) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(19286))))  severity failure;
	assert RAM(19287) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19287))))  severity failure;
	assert RAM(19288) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(19288))))  severity failure;
	assert RAM(19289) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19289))))  severity failure;
	assert RAM(19290) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(19290))))  severity failure;
	assert RAM(19291) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19291))))  severity failure;
	assert RAM(19292) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19292))))  severity failure;
	assert RAM(19293) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(19293))))  severity failure;
	assert RAM(19294) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(19294))))  severity failure;
	assert RAM(19295) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19295))))  severity failure;
	assert RAM(19296) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(19296))))  severity failure;
	assert RAM(19297) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19297))))  severity failure;
	assert RAM(19298) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19298))))  severity failure;
	assert RAM(19299) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(19299))))  severity failure;
	assert RAM(19300) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(19300))))  severity failure;
	assert RAM(19301) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(19301))))  severity failure;
	assert RAM(19302) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19302))))  severity failure;
	assert RAM(19303) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(19303))))  severity failure;
	assert RAM(19304) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19304))))  severity failure;
	assert RAM(19305) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19305))))  severity failure;
	assert RAM(19306) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(19306))))  severity failure;
	assert RAM(19307) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(19307))))  severity failure;
	assert RAM(19308) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(19308))))  severity failure;
	assert RAM(19309) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(19309))))  severity failure;
	assert RAM(19310) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(19310))))  severity failure;
	assert RAM(19311) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(19311))))  severity failure;
	assert RAM(19312) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19312))))  severity failure;
	assert RAM(19313) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(19313))))  severity failure;
	assert RAM(19314) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19314))))  severity failure;
	assert RAM(19315) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(19315))))  severity failure;
	assert RAM(19316) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(19316))))  severity failure;
	assert RAM(19317) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(19317))))  severity failure;
	assert RAM(19318) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(19318))))  severity failure;
	assert RAM(19319) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(19319))))  severity failure;
	assert RAM(19320) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19320))))  severity failure;
	assert RAM(19321) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(19321))))  severity failure;
	assert RAM(19322) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(19322))))  severity failure;
	assert RAM(19323) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(19323))))  severity failure;
	assert RAM(19324) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(19324))))  severity failure;
	assert RAM(19325) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(19325))))  severity failure;
	assert RAM(19326) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(19326))))  severity failure;
	assert RAM(19327) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(19327))))  severity failure;
	assert RAM(19328) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19328))))  severity failure;
	assert RAM(19329) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(19329))))  severity failure;
	assert RAM(19330) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(19330))))  severity failure;
	assert RAM(19331) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(19331))))  severity failure;
	assert RAM(19332) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(19332))))  severity failure;
	assert RAM(19333) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19333))))  severity failure;
	assert RAM(19334) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(19334))))  severity failure;
	assert RAM(19335) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19335))))  severity failure;
	assert RAM(19336) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(19336))))  severity failure;
	assert RAM(19337) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(19337))))  severity failure;
	assert RAM(19338) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19338))))  severity failure;
	assert RAM(19339) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(19339))))  severity failure;
	assert RAM(19340) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19340))))  severity failure;
	assert RAM(19341) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(19341))))  severity failure;
	assert RAM(19342) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19342))))  severity failure;
	assert RAM(19343) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19343))))  severity failure;
	assert RAM(19344) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19344))))  severity failure;
	assert RAM(19345) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19345))))  severity failure;
	assert RAM(19346) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(19346))))  severity failure;
	assert RAM(19347) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19347))))  severity failure;
	assert RAM(19348) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(19348))))  severity failure;
	assert RAM(19349) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19349))))  severity failure;
	assert RAM(19350) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(19350))))  severity failure;
	assert RAM(19351) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(19351))))  severity failure;
	assert RAM(19352) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(19352))))  severity failure;
	assert RAM(19353) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(19353))))  severity failure;
	assert RAM(19354) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(19354))))  severity failure;
	assert RAM(19355) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19355))))  severity failure;
	assert RAM(19356) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(19356))))  severity failure;
	assert RAM(19357) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(19357))))  severity failure;
	assert RAM(19358) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(19358))))  severity failure;
	assert RAM(19359) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(19359))))  severity failure;
	assert RAM(19360) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(19360))))  severity failure;
	assert RAM(19361) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(19361))))  severity failure;
	assert RAM(19362) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19362))))  severity failure;
	assert RAM(19363) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(19363))))  severity failure;
	assert RAM(19364) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(19364))))  severity failure;
	assert RAM(19365) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(19365))))  severity failure;
	assert RAM(19366) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(19366))))  severity failure;
	assert RAM(19367) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(19367))))  severity failure;
	assert RAM(19368) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(19368))))  severity failure;
	assert RAM(19369) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19369))))  severity failure;
	assert RAM(19370) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(19370))))  severity failure;
	assert RAM(19371) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19371))))  severity failure;
	assert RAM(19372) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(19372))))  severity failure;
	assert RAM(19373) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(19373))))  severity failure;
	assert RAM(19374) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(19374))))  severity failure;
	assert RAM(19375) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(19375))))  severity failure;
	assert RAM(19376) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(19376))))  severity failure;
	assert RAM(19377) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(19377))))  severity failure;
	assert RAM(19378) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(19378))))  severity failure;
	assert RAM(19379) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(19379))))  severity failure;
	assert RAM(19380) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(19380))))  severity failure;
	assert RAM(19381) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(19381))))  severity failure;
	assert RAM(19382) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(19382))))  severity failure;
	assert RAM(19383) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(19383))))  severity failure;
	assert RAM(19384) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19384))))  severity failure;
	assert RAM(19385) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(19385))))  severity failure;
	assert RAM(19386) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(19386))))  severity failure;
	assert RAM(19387) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(19387))))  severity failure;
	assert RAM(19388) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(19388))))  severity failure;
	assert RAM(19389) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(19389))))  severity failure;
	assert RAM(19390) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(19390))))  severity failure;
	assert RAM(19391) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19391))))  severity failure;
	assert RAM(19392) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19392))))  severity failure;
	assert RAM(19393) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(19393))))  severity failure;
	assert RAM(19394) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(19394))))  severity failure;
	assert RAM(19395) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(19395))))  severity failure;
	assert RAM(19396) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19396))))  severity failure;
	assert RAM(19397) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(19397))))  severity failure;
	assert RAM(19398) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(19398))))  severity failure;
	assert RAM(19399) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(19399))))  severity failure;
	assert RAM(19400) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(19400))))  severity failure;
	assert RAM(19401) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(19401))))  severity failure;
	assert RAM(19402) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(19402))))  severity failure;
	assert RAM(19403) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19403))))  severity failure;
	assert RAM(19404) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(19404))))  severity failure;
	assert RAM(19405) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19405))))  severity failure;
	assert RAM(19406) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19406))))  severity failure;
	assert RAM(19407) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(19407))))  severity failure;
	assert RAM(19408) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19408))))  severity failure;
	assert RAM(19409) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19409))))  severity failure;
	assert RAM(19410) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19410))))  severity failure;
	assert RAM(19411) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(19411))))  severity failure;
	assert RAM(19412) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(19412))))  severity failure;
	assert RAM(19413) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(19413))))  severity failure;
	assert RAM(19414) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(19414))))  severity failure;
	assert RAM(19415) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(19415))))  severity failure;
	assert RAM(19416) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(19416))))  severity failure;
	assert RAM(19417) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(19417))))  severity failure;
	assert RAM(19418) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19418))))  severity failure;
	assert RAM(19419) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(19419))))  severity failure;
	assert RAM(19420) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(19420))))  severity failure;
	assert RAM(19421) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(19421))))  severity failure;
	assert RAM(19422) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(19422))))  severity failure;
	assert RAM(19423) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(19423))))  severity failure;
	assert RAM(19424) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(19424))))  severity failure;
	assert RAM(19425) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(19425))))  severity failure;
	assert RAM(19426) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(19426))))  severity failure;
	assert RAM(19427) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(19427))))  severity failure;
	assert RAM(19428) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(19428))))  severity failure;
	assert RAM(19429) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19429))))  severity failure;
	assert RAM(19430) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(19430))))  severity failure;
	assert RAM(19431) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(19431))))  severity failure;
	assert RAM(19432) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19432))))  severity failure;
	assert RAM(19433) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(19433))))  severity failure;
	assert RAM(19434) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(19434))))  severity failure;
	assert RAM(19435) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(19435))))  severity failure;
	assert RAM(19436) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(19436))))  severity failure;
	assert RAM(19437) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19437))))  severity failure;
	assert RAM(19438) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(19438))))  severity failure;
	assert RAM(19439) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(19439))))  severity failure;
	assert RAM(19440) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(19440))))  severity failure;
	assert RAM(19441) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(19441))))  severity failure;
	assert RAM(19442) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(19442))))  severity failure;
	assert RAM(19443) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19443))))  severity failure;
	assert RAM(19444) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(19444))))  severity failure;
	assert RAM(19445) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19445))))  severity failure;
	assert RAM(19446) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(19446))))  severity failure;
	assert RAM(19447) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(19447))))  severity failure;
	assert RAM(19448) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(19448))))  severity failure;
	assert RAM(19449) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(19449))))  severity failure;
	assert RAM(19450) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(19450))))  severity failure;
	assert RAM(19451) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(19451))))  severity failure;
	assert RAM(19452) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19452))))  severity failure;
	assert RAM(19453) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(19453))))  severity failure;
	assert RAM(19454) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(19454))))  severity failure;
	assert RAM(19455) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(19455))))  severity failure;
	assert RAM(19456) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(19456))))  severity failure;
	assert RAM(19457) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(19457))))  severity failure;
	assert RAM(19458) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(19458))))  severity failure;
	assert RAM(19459) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(19459))))  severity failure;
	assert RAM(19460) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19460))))  severity failure;
	assert RAM(19461) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(19461))))  severity failure;
	assert RAM(19462) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(19462))))  severity failure;
	assert RAM(19463) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(19463))))  severity failure;
	assert RAM(19464) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(19464))))  severity failure;
	assert RAM(19465) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(19465))))  severity failure;
	assert RAM(19466) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19466))))  severity failure;
	assert RAM(19467) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(19467))))  severity failure;
	assert RAM(19468) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(19468))))  severity failure;
	assert RAM(19469) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(19469))))  severity failure;
	assert RAM(19470) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19470))))  severity failure;
	assert RAM(19471) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(19471))))  severity failure;
	assert RAM(19472) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(19472))))  severity failure;
	assert RAM(19473) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(19473))))  severity failure;
	assert RAM(19474) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19474))))  severity failure;
	assert RAM(19475) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(19475))))  severity failure;
	assert RAM(19476) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19476))))  severity failure;
	assert RAM(19477) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(19477))))  severity failure;
	assert RAM(19478) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(19478))))  severity failure;
	assert RAM(19479) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(19479))))  severity failure;
	assert RAM(19480) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19480))))  severity failure;
	assert RAM(19481) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(19481))))  severity failure;
	assert RAM(19482) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19482))))  severity failure;
	assert RAM(19483) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(19483))))  severity failure;
	assert RAM(19484) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19484))))  severity failure;
	assert RAM(19485) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(19485))))  severity failure;
	assert RAM(19486) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(19486))))  severity failure;
	assert RAM(19487) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(19487))))  severity failure;
	assert RAM(19488) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19488))))  severity failure;
	assert RAM(19489) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(19489))))  severity failure;
	assert RAM(19490) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(19490))))  severity failure;
	assert RAM(19491) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19491))))  severity failure;
	assert RAM(19492) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(19492))))  severity failure;
	assert RAM(19493) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(19493))))  severity failure;
	assert RAM(19494) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(19494))))  severity failure;
	assert RAM(19495) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19495))))  severity failure;
	assert RAM(19496) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(19496))))  severity failure;
	assert RAM(19497) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(19497))))  severity failure;
	assert RAM(19498) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(19498))))  severity failure;
	assert RAM(19499) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(19499))))  severity failure;
	assert RAM(19500) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(19500))))  severity failure;
	assert RAM(19501) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(19501))))  severity failure;
	assert RAM(19502) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19502))))  severity failure;
	assert RAM(19503) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(19503))))  severity failure;
	assert RAM(19504) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19504))))  severity failure;
	assert RAM(19505) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(19505))))  severity failure;
	assert RAM(19506) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(19506))))  severity failure;
	assert RAM(19507) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19507))))  severity failure;
	assert RAM(19508) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(19508))))  severity failure;
	assert RAM(19509) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(19509))))  severity failure;
	assert RAM(19510) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(19510))))  severity failure;
	assert RAM(19511) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(19511))))  severity failure;
	assert RAM(19512) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(19512))))  severity failure;
	assert RAM(19513) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(19513))))  severity failure;
	assert RAM(19514) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(19514))))  severity failure;
	assert RAM(19515) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19515))))  severity failure;
	assert RAM(19516) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(19516))))  severity failure;
	assert RAM(19517) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19517))))  severity failure;
	assert RAM(19518) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19518))))  severity failure;
	assert RAM(19519) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(19519))))  severity failure;
	assert RAM(19520) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(19520))))  severity failure;
	assert RAM(19521) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19521))))  severity failure;
	assert RAM(19522) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(19522))))  severity failure;
	assert RAM(19523) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(19523))))  severity failure;
	assert RAM(19524) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(19524))))  severity failure;
	assert RAM(19525) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(19525))))  severity failure;
	assert RAM(19526) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(19526))))  severity failure;
	assert RAM(19527) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(19527))))  severity failure;
	assert RAM(19528) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(19528))))  severity failure;
	assert RAM(19529) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(19529))))  severity failure;
	assert RAM(19530) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(19530))))  severity failure;
	assert RAM(19531) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19531))))  severity failure;
	assert RAM(19532) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(19532))))  severity failure;
	assert RAM(19533) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(19533))))  severity failure;
	assert RAM(19534) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19534))))  severity failure;
	assert RAM(19535) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(19535))))  severity failure;
	assert RAM(19536) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(19536))))  severity failure;
	assert RAM(19537) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(19537))))  severity failure;
	assert RAM(19538) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(19538))))  severity failure;
	assert RAM(19539) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19539))))  severity failure;
	assert RAM(19540) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(19540))))  severity failure;
	assert RAM(19541) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(19541))))  severity failure;
	assert RAM(19542) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(19542))))  severity failure;
	assert RAM(19543) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(19543))))  severity failure;
	assert RAM(19544) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19544))))  severity failure;
	assert RAM(19545) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(19545))))  severity failure;
	assert RAM(19546) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19546))))  severity failure;
	assert RAM(19547) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(19547))))  severity failure;
	assert RAM(19548) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19548))))  severity failure;
	assert RAM(19549) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(19549))))  severity failure;
	assert RAM(19550) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(19550))))  severity failure;
	assert RAM(19551) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(19551))))  severity failure;
	assert RAM(19552) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(19552))))  severity failure;
	assert RAM(19553) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(19553))))  severity failure;
	assert RAM(19554) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(19554))))  severity failure;
	assert RAM(19555) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(19555))))  severity failure;
	assert RAM(19556) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(19556))))  severity failure;
	assert RAM(19557) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(19557))))  severity failure;
	assert RAM(19558) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(19558))))  severity failure;
	assert RAM(19559) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(19559))))  severity failure;
	assert RAM(19560) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(19560))))  severity failure;
	assert RAM(19561) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(19561))))  severity failure;
	assert RAM(19562) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(19562))))  severity failure;
	assert RAM(19563) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(19563))))  severity failure;
	assert RAM(19564) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(19564))))  severity failure;
	assert RAM(19565) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(19565))))  severity failure;
	assert RAM(19566) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19566))))  severity failure;
	assert RAM(19567) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(19567))))  severity failure;
	assert RAM(19568) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(19568))))  severity failure;
	assert RAM(19569) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(19569))))  severity failure;
	assert RAM(19570) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(19570))))  severity failure;
	assert RAM(19571) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(19571))))  severity failure;
	assert RAM(19572) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(19572))))  severity failure;
	assert RAM(19573) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19573))))  severity failure;
	assert RAM(19574) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(19574))))  severity failure;
	assert RAM(19575) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(19575))))  severity failure;
	assert RAM(19576) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(19576))))  severity failure;
	assert RAM(19577) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19577))))  severity failure;
	assert RAM(19578) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(19578))))  severity failure;
	assert RAM(19579) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(19579))))  severity failure;
	assert RAM(19580) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(19580))))  severity failure;
	assert RAM(19581) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19581))))  severity failure;
	assert RAM(19582) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(19582))))  severity failure;
	assert RAM(19583) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(19583))))  severity failure;
	assert RAM(19584) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19584))))  severity failure;
	assert RAM(19585) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19585))))  severity failure;
	assert RAM(19586) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(19586))))  severity failure;
	assert RAM(19587) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(19587))))  severity failure;
	assert RAM(19588) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19588))))  severity failure;
	assert RAM(19589) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(19589))))  severity failure;
	assert RAM(19590) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(19590))))  severity failure;
	assert RAM(19591) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(19591))))  severity failure;
	assert RAM(19592) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19592))))  severity failure;
	assert RAM(19593) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(19593))))  severity failure;
	assert RAM(19594) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(19594))))  severity failure;
	assert RAM(19595) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(19595))))  severity failure;
	assert RAM(19596) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(19596))))  severity failure;
	assert RAM(19597) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19597))))  severity failure;
	assert RAM(19598) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(19598))))  severity failure;
	assert RAM(19599) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19599))))  severity failure;
	assert RAM(19600) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(19600))))  severity failure;
	assert RAM(19601) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(19601))))  severity failure;
	assert RAM(19602) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(19602))))  severity failure;
	assert RAM(19603) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(19603))))  severity failure;
	assert RAM(19604) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(19604))))  severity failure;
	assert RAM(19605) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(19605))))  severity failure;
	assert RAM(19606) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(19606))))  severity failure;
	assert RAM(19607) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19607))))  severity failure;
	assert RAM(19608) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(19608))))  severity failure;
	assert RAM(19609) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(19609))))  severity failure;
	assert RAM(19610) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19610))))  severity failure;
	assert RAM(19611) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(19611))))  severity failure;
	assert RAM(19612) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19612))))  severity failure;
	assert RAM(19613) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(19613))))  severity failure;
	assert RAM(19614) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(19614))))  severity failure;
	assert RAM(19615) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(19615))))  severity failure;
	assert RAM(19616) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19616))))  severity failure;
	assert RAM(19617) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(19617))))  severity failure;
	assert RAM(19618) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(19618))))  severity failure;
	assert RAM(19619) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19619))))  severity failure;
	assert RAM(19620) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(19620))))  severity failure;
	assert RAM(19621) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(19621))))  severity failure;
	assert RAM(19622) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19622))))  severity failure;
	assert RAM(19623) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19623))))  severity failure;
	assert RAM(19624) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(19624))))  severity failure;
	assert RAM(19625) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(19625))))  severity failure;
	assert RAM(19626) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(19626))))  severity failure;
	assert RAM(19627) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(19627))))  severity failure;
	assert RAM(19628) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19628))))  severity failure;
	assert RAM(19629) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(19629))))  severity failure;
	assert RAM(19630) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(19630))))  severity failure;
	assert RAM(19631) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(19631))))  severity failure;
	assert RAM(19632) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(19632))))  severity failure;
	assert RAM(19633) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(19633))))  severity failure;
	assert RAM(19634) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(19634))))  severity failure;
	assert RAM(19635) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(19635))))  severity failure;
	assert RAM(19636) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(19636))))  severity failure;
	assert RAM(19637) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(19637))))  severity failure;
	assert RAM(19638) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(19638))))  severity failure;
	assert RAM(19639) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(19639))))  severity failure;
	assert RAM(19640) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(19640))))  severity failure;
	assert RAM(19641) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(19641))))  severity failure;
	assert RAM(19642) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19642))))  severity failure;
	assert RAM(19643) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(19643))))  severity failure;
	assert RAM(19644) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19644))))  severity failure;
	assert RAM(19645) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(19645))))  severity failure;
	assert RAM(19646) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(19646))))  severity failure;
	assert RAM(19647) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19647))))  severity failure;
	assert RAM(19648) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(19648))))  severity failure;
	assert RAM(19649) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(19649))))  severity failure;
	assert RAM(19650) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19650))))  severity failure;
	assert RAM(19651) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(19651))))  severity failure;
	assert RAM(19652) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19652))))  severity failure;
	assert RAM(19653) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(19653))))  severity failure;
	assert RAM(19654) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(19654))))  severity failure;
	assert RAM(19655) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(19655))))  severity failure;
	assert RAM(19656) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(19656))))  severity failure;
	assert RAM(19657) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(19657))))  severity failure;
	assert RAM(19658) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(19658))))  severity failure;
	assert RAM(19659) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19659))))  severity failure;
	assert RAM(19660) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(19660))))  severity failure;
	assert RAM(19661) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(19661))))  severity failure;
	assert RAM(19662) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(19662))))  severity failure;
	assert RAM(19663) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(19663))))  severity failure;
	assert RAM(19664) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(19664))))  severity failure;
	assert RAM(19665) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(19665))))  severity failure;
	assert RAM(19666) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(19666))))  severity failure;
	assert RAM(19667) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(19667))))  severity failure;
	assert RAM(19668) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(19668))))  severity failure;
	assert RAM(19669) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(19669))))  severity failure;
	assert RAM(19670) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(19670))))  severity failure;
	assert RAM(19671) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(19671))))  severity failure;
	assert RAM(19672) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(19672))))  severity failure;
	assert RAM(19673) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(19673))))  severity failure;
	assert RAM(19674) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(19674))))  severity failure;
	assert RAM(19675) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(19675))))  severity failure;
	assert RAM(19676) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(19676))))  severity failure;
	assert RAM(19677) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19677))))  severity failure;
	assert RAM(19678) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(19678))))  severity failure;
	assert RAM(19679) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19679))))  severity failure;
	assert RAM(19680) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(19680))))  severity failure;
	assert RAM(19681) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(19681))))  severity failure;
	assert RAM(19682) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(19682))))  severity failure;
	assert RAM(19683) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(19683))))  severity failure;
	assert RAM(19684) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(19684))))  severity failure;
	assert RAM(19685) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(19685))))  severity failure;
	assert RAM(19686) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19686))))  severity failure;
	assert RAM(19687) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(19687))))  severity failure;
	assert RAM(19688) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19688))))  severity failure;
	assert RAM(19689) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(19689))))  severity failure;
	assert RAM(19690) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(19690))))  severity failure;
	assert RAM(19691) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19691))))  severity failure;
	assert RAM(19692) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(19692))))  severity failure;
	assert RAM(19693) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19693))))  severity failure;
	assert RAM(19694) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(19694))))  severity failure;
	assert RAM(19695) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(19695))))  severity failure;
	assert RAM(19696) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(19696))))  severity failure;
	assert RAM(19697) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(19697))))  severity failure;
	assert RAM(19698) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(19698))))  severity failure;
	assert RAM(19699) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(19699))))  severity failure;
	assert RAM(19700) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(19700))))  severity failure;
	assert RAM(19701) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(19701))))  severity failure;
	assert RAM(19702) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19702))))  severity failure;
	assert RAM(19703) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(19703))))  severity failure;
	assert RAM(19704) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(19704))))  severity failure;
	assert RAM(19705) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(19705))))  severity failure;
	assert RAM(19706) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(19706))))  severity failure;
	assert RAM(19707) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(19707))))  severity failure;
	assert RAM(19708) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(19708))))  severity failure;
	assert RAM(19709) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(19709))))  severity failure;
	assert RAM(19710) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(19710))))  severity failure;
	assert RAM(19711) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(19711))))  severity failure;
	assert RAM(19712) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(19712))))  severity failure;
	assert RAM(19713) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(19713))))  severity failure;
	assert RAM(19714) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(19714))))  severity failure;
	assert RAM(19715) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(19715))))  severity failure;
	assert RAM(19716) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(19716))))  severity failure;
	assert RAM(19717) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(19717))))  severity failure;
	assert RAM(19718) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(19718))))  severity failure;
	assert RAM(19719) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(19719))))  severity failure;
	assert RAM(19720) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(19720))))  severity failure;
	assert RAM(19721) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(19721))))  severity failure;
	assert RAM(19722) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(19722))))  severity failure;
	assert RAM(19723) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(19723))))  severity failure;
	assert RAM(19724) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(19724))))  severity failure;
	assert RAM(19725) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(19725))))  severity failure;
	assert RAM(19726) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(19726))))  severity failure;
	assert RAM(19727) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19727))))  severity failure;
	assert RAM(19728) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(19728))))  severity failure;
	assert RAM(19729) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19729))))  severity failure;
	assert RAM(19730) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19730))))  severity failure;
	assert RAM(19731) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(19731))))  severity failure;
	assert RAM(19732) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(19732))))  severity failure;
	assert RAM(19733) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(19733))))  severity failure;
	assert RAM(19734) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(19734))))  severity failure;
	assert RAM(19735) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(19735))))  severity failure;
	assert RAM(19736) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(19736))))  severity failure;
	assert RAM(19737) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(19737))))  severity failure;
	assert RAM(19738) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(19738))))  severity failure;
	assert RAM(19739) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(19739))))  severity failure;
	assert RAM(19740) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(19740))))  severity failure;
	assert RAM(19741) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(19741))))  severity failure;
	assert RAM(19742) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(19742))))  severity failure;
	assert RAM(19743) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(19743))))  severity failure;
	assert RAM(19744) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19744))))  severity failure;
	assert RAM(19745) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(19745))))  severity failure;
	assert RAM(19746) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19746))))  severity failure;
	assert RAM(19747) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(19747))))  severity failure;
	assert RAM(19748) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(19748))))  severity failure;
	assert RAM(19749) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(19749))))  severity failure;
	assert RAM(19750) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(19750))))  severity failure;
	assert RAM(19751) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(19751))))  severity failure;
	assert RAM(19752) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(19752))))  severity failure;
	assert RAM(19753) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19753))))  severity failure;
	assert RAM(19754) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(19754))))  severity failure;
	assert RAM(19755) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(19755))))  severity failure;
	assert RAM(19756) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(19756))))  severity failure;
	assert RAM(19757) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19757))))  severity failure;
	assert RAM(19758) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(19758))))  severity failure;
	assert RAM(19759) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(19759))))  severity failure;
	assert RAM(19760) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(19760))))  severity failure;
	assert RAM(19761) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(19761))))  severity failure;
	assert RAM(19762) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(19762))))  severity failure;
	assert RAM(19763) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19763))))  severity failure;
	assert RAM(19764) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(19764))))  severity failure;
	assert RAM(19765) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(19765))))  severity failure;
	assert RAM(19766) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(19766))))  severity failure;
	assert RAM(19767) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(19767))))  severity failure;
	assert RAM(19768) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19768))))  severity failure;
	assert RAM(19769) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(19769))))  severity failure;
	assert RAM(19770) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(19770))))  severity failure;
	assert RAM(19771) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(19771))))  severity failure;
	assert RAM(19772) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(19772))))  severity failure;
	assert RAM(19773) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(19773))))  severity failure;
	assert RAM(19774) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19774))))  severity failure;
	assert RAM(19775) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(19775))))  severity failure;
	assert RAM(19776) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(19776))))  severity failure;
	assert RAM(19777) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(19777))))  severity failure;
	assert RAM(19778) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19778))))  severity failure;
	assert RAM(19779) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(19779))))  severity failure;
	assert RAM(19780) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19780))))  severity failure;
	assert RAM(19781) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(19781))))  severity failure;
	assert RAM(19782) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19782))))  severity failure;
	assert RAM(19783) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(19783))))  severity failure;
	assert RAM(19784) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(19784))))  severity failure;
	assert RAM(19785) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(19785))))  severity failure;
	assert RAM(19786) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19786))))  severity failure;
	assert RAM(19787) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(19787))))  severity failure;
	assert RAM(19788) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(19788))))  severity failure;
	assert RAM(19789) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(19789))))  severity failure;
	assert RAM(19790) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19790))))  severity failure;
	assert RAM(19791) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(19791))))  severity failure;
	assert RAM(19792) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(19792))))  severity failure;
	assert RAM(19793) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(19793))))  severity failure;
	assert RAM(19794) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19794))))  severity failure;
	assert RAM(19795) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(19795))))  severity failure;
	assert RAM(19796) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(19796))))  severity failure;
	assert RAM(19797) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(19797))))  severity failure;
	assert RAM(19798) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(19798))))  severity failure;
	assert RAM(19799) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(19799))))  severity failure;
	assert RAM(19800) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(19800))))  severity failure;
	assert RAM(19801) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19801))))  severity failure;
	assert RAM(19802) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(19802))))  severity failure;
	assert RAM(19803) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(19803))))  severity failure;
	assert RAM(19804) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19804))))  severity failure;
	assert RAM(19805) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(19805))))  severity failure;
	assert RAM(19806) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(19806))))  severity failure;
	assert RAM(19807) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(19807))))  severity failure;
	assert RAM(19808) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(19808))))  severity failure;
	assert RAM(19809) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(19809))))  severity failure;
	assert RAM(19810) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(19810))))  severity failure;
	assert RAM(19811) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(19811))))  severity failure;
	assert RAM(19812) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(19812))))  severity failure;
	assert RAM(19813) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(19813))))  severity failure;
	assert RAM(19814) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(19814))))  severity failure;
	assert RAM(19815) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(19815))))  severity failure;
	assert RAM(19816) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19816))))  severity failure;
	assert RAM(19817) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(19817))))  severity failure;
	assert RAM(19818) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(19818))))  severity failure;
	assert RAM(19819) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(19819))))  severity failure;
	assert RAM(19820) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19820))))  severity failure;
	assert RAM(19821) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(19821))))  severity failure;
	assert RAM(19822) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(19822))))  severity failure;
	assert RAM(19823) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(19823))))  severity failure;
	assert RAM(19824) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(19824))))  severity failure;
	assert RAM(19825) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(19825))))  severity failure;
	assert RAM(19826) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(19826))))  severity failure;
	assert RAM(19827) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(19827))))  severity failure;
	assert RAM(19828) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(19828))))  severity failure;
	assert RAM(19829) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(19829))))  severity failure;
	assert RAM(19830) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(19830))))  severity failure;
	assert RAM(19831) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(19831))))  severity failure;
	assert RAM(19832) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(19832))))  severity failure;
	assert RAM(19833) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19833))))  severity failure;
	assert RAM(19834) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(19834))))  severity failure;
	assert RAM(19835) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(19835))))  severity failure;
	assert RAM(19836) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(19836))))  severity failure;
	assert RAM(19837) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19837))))  severity failure;
	assert RAM(19838) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(19838))))  severity failure;
	assert RAM(19839) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(19839))))  severity failure;
	assert RAM(19840) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(19840))))  severity failure;
	assert RAM(19841) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(19841))))  severity failure;
	assert RAM(19842) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(19842))))  severity failure;
	assert RAM(19843) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(19843))))  severity failure;
	assert RAM(19844) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(19844))))  severity failure;
	assert RAM(19845) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(19845))))  severity failure;
	assert RAM(19846) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19846))))  severity failure;
	assert RAM(19847) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19847))))  severity failure;
	assert RAM(19848) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(19848))))  severity failure;
	assert RAM(19849) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(19849))))  severity failure;
	assert RAM(19850) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(19850))))  severity failure;
	assert RAM(19851) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(19851))))  severity failure;
	assert RAM(19852) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(19852))))  severity failure;
	assert RAM(19853) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19853))))  severity failure;
	assert RAM(19854) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19854))))  severity failure;
	assert RAM(19855) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(19855))))  severity failure;
	assert RAM(19856) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(19856))))  severity failure;
	assert RAM(19857) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(19857))))  severity failure;
	assert RAM(19858) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19858))))  severity failure;
	assert RAM(19859) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(19859))))  severity failure;
	assert RAM(19860) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(19860))))  severity failure;
	assert RAM(19861) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(19861))))  severity failure;
	assert RAM(19862) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(19862))))  severity failure;
	assert RAM(19863) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(19863))))  severity failure;
	assert RAM(19864) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19864))))  severity failure;
	assert RAM(19865) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19865))))  severity failure;
	assert RAM(19866) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(19866))))  severity failure;
	assert RAM(19867) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(19867))))  severity failure;
	assert RAM(19868) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(19868))))  severity failure;
	assert RAM(19869) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19869))))  severity failure;
	assert RAM(19870) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19870))))  severity failure;
	assert RAM(19871) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(19871))))  severity failure;
	assert RAM(19872) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19872))))  severity failure;
	assert RAM(19873) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(19873))))  severity failure;
	assert RAM(19874) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(19874))))  severity failure;
	assert RAM(19875) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(19875))))  severity failure;
	assert RAM(19876) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(19876))))  severity failure;
	assert RAM(19877) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(19877))))  severity failure;
	assert RAM(19878) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(19878))))  severity failure;
	assert RAM(19879) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(19879))))  severity failure;
	assert RAM(19880) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(19880))))  severity failure;
	assert RAM(19881) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(19881))))  severity failure;
	assert RAM(19882) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(19882))))  severity failure;
	assert RAM(19883) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(19883))))  severity failure;
	assert RAM(19884) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(19884))))  severity failure;
	assert RAM(19885) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19885))))  severity failure;
	assert RAM(19886) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(19886))))  severity failure;
	assert RAM(19887) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(19887))))  severity failure;
	assert RAM(19888) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(19888))))  severity failure;
	assert RAM(19889) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(19889))))  severity failure;
	assert RAM(19890) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(19890))))  severity failure;
	assert RAM(19891) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19891))))  severity failure;
	assert RAM(19892) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(19892))))  severity failure;
	assert RAM(19893) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(19893))))  severity failure;
	assert RAM(19894) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(19894))))  severity failure;
	assert RAM(19895) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(19895))))  severity failure;
	assert RAM(19896) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(19896))))  severity failure;
	assert RAM(19897) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(19897))))  severity failure;
	assert RAM(19898) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(19898))))  severity failure;
	assert RAM(19899) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(19899))))  severity failure;
	assert RAM(19900) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(19900))))  severity failure;
	assert RAM(19901) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(19901))))  severity failure;
	assert RAM(19902) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19902))))  severity failure;
	assert RAM(19903) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(19903))))  severity failure;
	assert RAM(19904) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(19904))))  severity failure;
	assert RAM(19905) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(19905))))  severity failure;
	assert RAM(19906) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(19906))))  severity failure;
	assert RAM(19907) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(19907))))  severity failure;
	assert RAM(19908) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(19908))))  severity failure;
	assert RAM(19909) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(19909))))  severity failure;
	assert RAM(19910) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(19910))))  severity failure;
	assert RAM(19911) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(19911))))  severity failure;
	assert RAM(19912) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(19912))))  severity failure;
	assert RAM(19913) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(19913))))  severity failure;
	assert RAM(19914) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(19914))))  severity failure;
	assert RAM(19915) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(19915))))  severity failure;
	assert RAM(19916) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(19916))))  severity failure;
	assert RAM(19917) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(19917))))  severity failure;
	assert RAM(19918) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(19918))))  severity failure;
	assert RAM(19919) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19919))))  severity failure;
	assert RAM(19920) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(19920))))  severity failure;
	assert RAM(19921) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(19921))))  severity failure;
	assert RAM(19922) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19922))))  severity failure;
	assert RAM(19923) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(19923))))  severity failure;
	assert RAM(19924) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(19924))))  severity failure;
	assert RAM(19925) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(19925))))  severity failure;
	assert RAM(19926) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(19926))))  severity failure;
	assert RAM(19927) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(19927))))  severity failure;
	assert RAM(19928) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(19928))))  severity failure;
	assert RAM(19929) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(19929))))  severity failure;
	assert RAM(19930) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(19930))))  severity failure;
	assert RAM(19931) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(19931))))  severity failure;
	assert RAM(19932) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(19932))))  severity failure;
	assert RAM(19933) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(19933))))  severity failure;
	assert RAM(19934) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(19934))))  severity failure;
	assert RAM(19935) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(19935))))  severity failure;
	assert RAM(19936) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(19936))))  severity failure;
	assert RAM(19937) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(19937))))  severity failure;
	assert RAM(19938) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(19938))))  severity failure;
	assert RAM(19939) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19939))))  severity failure;
	assert RAM(19940) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(19940))))  severity failure;
	assert RAM(19941) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(19941))))  severity failure;
	assert RAM(19942) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19942))))  severity failure;
	assert RAM(19943) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(19943))))  severity failure;
	assert RAM(19944) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(19944))))  severity failure;
	assert RAM(19945) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19945))))  severity failure;
	assert RAM(19946) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(19946))))  severity failure;
	assert RAM(19947) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(19947))))  severity failure;
	assert RAM(19948) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(19948))))  severity failure;
	assert RAM(19949) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(19949))))  severity failure;
	assert RAM(19950) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(19950))))  severity failure;
	assert RAM(19951) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(19951))))  severity failure;
	assert RAM(19952) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(19952))))  severity failure;
	assert RAM(19953) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(19953))))  severity failure;
	assert RAM(19954) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(19954))))  severity failure;
	assert RAM(19955) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(19955))))  severity failure;
	assert RAM(19956) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(19956))))  severity failure;
	assert RAM(19957) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(19957))))  severity failure;
	assert RAM(19958) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(19958))))  severity failure;
	assert RAM(19959) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(19959))))  severity failure;
	assert RAM(19960) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(19960))))  severity failure;
	assert RAM(19961) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(19961))))  severity failure;
	assert RAM(19962) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(19962))))  severity failure;
	assert RAM(19963) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(19963))))  severity failure;
	assert RAM(19964) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(19964))))  severity failure;
	assert RAM(19965) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(19965))))  severity failure;
	assert RAM(19966) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(19966))))  severity failure;
	assert RAM(19967) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(19967))))  severity failure;
	assert RAM(19968) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(19968))))  severity failure;
	assert RAM(19969) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(19969))))  severity failure;
	assert RAM(19970) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(19970))))  severity failure;
	assert RAM(19971) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(19971))))  severity failure;
	assert RAM(19972) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(19972))))  severity failure;
	assert RAM(19973) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(19973))))  severity failure;
	assert RAM(19974) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(19974))))  severity failure;
	assert RAM(19975) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(19975))))  severity failure;
	assert RAM(19976) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(19976))))  severity failure;
	assert RAM(19977) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(19977))))  severity failure;
	assert RAM(19978) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(19978))))  severity failure;
	assert RAM(19979) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(19979))))  severity failure;
	assert RAM(19980) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(19980))))  severity failure;
	assert RAM(19981) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(19981))))  severity failure;
	assert RAM(19982) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(19982))))  severity failure;
	assert RAM(19983) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(19983))))  severity failure;
	assert RAM(19984) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(19984))))  severity failure;
	assert RAM(19985) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(19985))))  severity failure;
	assert RAM(19986) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(19986))))  severity failure;
	assert RAM(19987) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(19987))))  severity failure;
	assert RAM(19988) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(19988))))  severity failure;
	assert RAM(19989) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(19989))))  severity failure;
	assert RAM(19990) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(19990))))  severity failure;
	assert RAM(19991) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(19991))))  severity failure;
	assert RAM(19992) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(19992))))  severity failure;
	assert RAM(19993) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(19993))))  severity failure;
	assert RAM(19994) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(19994))))  severity failure;
	assert RAM(19995) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(19995))))  severity failure;
	assert RAM(19996) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(19996))))  severity failure;
	assert RAM(19997) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(19997))))  severity failure;
	assert RAM(19998) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(19998))))  severity failure;
	assert RAM(19999) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(19999))))  severity failure;
	assert RAM(20000) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(20000))))  severity failure;
	assert RAM(20001) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(20001))))  severity failure;
	assert RAM(20002) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(20002))))  severity failure;
	assert RAM(20003) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20003))))  severity failure;
	assert RAM(20004) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(20004))))  severity failure;
	assert RAM(20005) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(20005))))  severity failure;
	assert RAM(20006) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20006))))  severity failure;
	assert RAM(20007) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(20007))))  severity failure;
	assert RAM(20008) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(20008))))  severity failure;
	assert RAM(20009) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20009))))  severity failure;
	assert RAM(20010) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(20010))))  severity failure;
	assert RAM(20011) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(20011))))  severity failure;
	assert RAM(20012) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20012))))  severity failure;
	assert RAM(20013) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(20013))))  severity failure;
	assert RAM(20014) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(20014))))  severity failure;
	assert RAM(20015) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20015))))  severity failure;
	assert RAM(20016) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(20016))))  severity failure;
	assert RAM(20017) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(20017))))  severity failure;
	assert RAM(20018) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(20018))))  severity failure;
	assert RAM(20019) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(20019))))  severity failure;
	assert RAM(20020) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(20020))))  severity failure;
	assert RAM(20021) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(20021))))  severity failure;
	assert RAM(20022) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20022))))  severity failure;
	assert RAM(20023) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(20023))))  severity failure;
	assert RAM(20024) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20024))))  severity failure;
	assert RAM(20025) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(20025))))  severity failure;
	assert RAM(20026) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(20026))))  severity failure;
	assert RAM(20027) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(20027))))  severity failure;
	assert RAM(20028) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20028))))  severity failure;
	assert RAM(20029) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20029))))  severity failure;
	assert RAM(20030) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20030))))  severity failure;
	assert RAM(20031) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(20031))))  severity failure;
	assert RAM(20032) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(20032))))  severity failure;
	assert RAM(20033) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20033))))  severity failure;
	assert RAM(20034) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(20034))))  severity failure;
	assert RAM(20035) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20035))))  severity failure;
	assert RAM(20036) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(20036))))  severity failure;
	assert RAM(20037) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(20037))))  severity failure;
	assert RAM(20038) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(20038))))  severity failure;
	assert RAM(20039) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20039))))  severity failure;
	assert RAM(20040) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(20040))))  severity failure;
	assert RAM(20041) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(20041))))  severity failure;
	assert RAM(20042) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20042))))  severity failure;
	assert RAM(20043) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(20043))))  severity failure;
	assert RAM(20044) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20044))))  severity failure;
	assert RAM(20045) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20045))))  severity failure;
	assert RAM(20046) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20046))))  severity failure;
	assert RAM(20047) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(20047))))  severity failure;
	assert RAM(20048) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20048))))  severity failure;
	assert RAM(20049) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(20049))))  severity failure;
	assert RAM(20050) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(20050))))  severity failure;
	assert RAM(20051) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(20051))))  severity failure;
	assert RAM(20052) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(20052))))  severity failure;
	assert RAM(20053) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(20053))))  severity failure;
	assert RAM(20054) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(20054))))  severity failure;
	assert RAM(20055) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(20055))))  severity failure;
	assert RAM(20056) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(20056))))  severity failure;
	assert RAM(20057) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(20057))))  severity failure;
	assert RAM(20058) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(20058))))  severity failure;
	assert RAM(20059) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(20059))))  severity failure;
	assert RAM(20060) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(20060))))  severity failure;
	assert RAM(20061) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(20061))))  severity failure;
	assert RAM(20062) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(20062))))  severity failure;
	assert RAM(20063) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(20063))))  severity failure;
	assert RAM(20064) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(20064))))  severity failure;
	assert RAM(20065) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(20065))))  severity failure;
	assert RAM(20066) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20066))))  severity failure;
	assert RAM(20067) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(20067))))  severity failure;
	assert RAM(20068) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20068))))  severity failure;
	assert RAM(20069) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(20069))))  severity failure;
	assert RAM(20070) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20070))))  severity failure;
	assert RAM(20071) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(20071))))  severity failure;
	assert RAM(20072) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(20072))))  severity failure;
	assert RAM(20073) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(20073))))  severity failure;
	assert RAM(20074) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(20074))))  severity failure;
	assert RAM(20075) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(20075))))  severity failure;
	assert RAM(20076) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(20076))))  severity failure;
	assert RAM(20077) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(20077))))  severity failure;
	assert RAM(20078) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(20078))))  severity failure;
	assert RAM(20079) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(20079))))  severity failure;
	assert RAM(20080) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20080))))  severity failure;
	assert RAM(20081) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(20081))))  severity failure;
	assert RAM(20082) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(20082))))  severity failure;
	assert RAM(20083) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(20083))))  severity failure;
	assert RAM(20084) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(20084))))  severity failure;
	assert RAM(20085) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(20085))))  severity failure;
	assert RAM(20086) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(20086))))  severity failure;
	assert RAM(20087) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(20087))))  severity failure;
	assert RAM(20088) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20088))))  severity failure;
	assert RAM(20089) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(20089))))  severity failure;
	assert RAM(20090) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(20090))))  severity failure;
	assert RAM(20091) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(20091))))  severity failure;
	assert RAM(20092) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(20092))))  severity failure;
	assert RAM(20093) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20093))))  severity failure;
	assert RAM(20094) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(20094))))  severity failure;
	assert RAM(20095) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(20095))))  severity failure;
	assert RAM(20096) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(20096))))  severity failure;
	assert RAM(20097) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(20097))))  severity failure;
	assert RAM(20098) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20098))))  severity failure;
	assert RAM(20099) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(20099))))  severity failure;
	assert RAM(20100) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(20100))))  severity failure;
	assert RAM(20101) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(20101))))  severity failure;
	assert RAM(20102) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20102))))  severity failure;
	assert RAM(20103) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20103))))  severity failure;
	assert RAM(20104) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(20104))))  severity failure;
	assert RAM(20105) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(20105))))  severity failure;
	assert RAM(20106) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(20106))))  severity failure;
	assert RAM(20107) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(20107))))  severity failure;
	assert RAM(20108) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(20108))))  severity failure;
	assert RAM(20109) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20109))))  severity failure;
	assert RAM(20110) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20110))))  severity failure;
	assert RAM(20111) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(20111))))  severity failure;
	assert RAM(20112) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(20112))))  severity failure;
	assert RAM(20113) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(20113))))  severity failure;
	assert RAM(20114) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(20114))))  severity failure;
	assert RAM(20115) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(20115))))  severity failure;
	assert RAM(20116) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(20116))))  severity failure;
	assert RAM(20117) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(20117))))  severity failure;
	assert RAM(20118) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(20118))))  severity failure;
	assert RAM(20119) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20119))))  severity failure;
	assert RAM(20120) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(20120))))  severity failure;
	assert RAM(20121) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(20121))))  severity failure;
	assert RAM(20122) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(20122))))  severity failure;
	assert RAM(20123) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(20123))))  severity failure;
	assert RAM(20124) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(20124))))  severity failure;
	assert RAM(20125) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(20125))))  severity failure;
	assert RAM(20126) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20126))))  severity failure;
	assert RAM(20127) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20127))))  severity failure;
	assert RAM(20128) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(20128))))  severity failure;
	assert RAM(20129) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20129))))  severity failure;
	assert RAM(20130) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20130))))  severity failure;
	assert RAM(20131) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(20131))))  severity failure;
	assert RAM(20132) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(20132))))  severity failure;
	assert RAM(20133) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(20133))))  severity failure;
	assert RAM(20134) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(20134))))  severity failure;
	assert RAM(20135) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(20135))))  severity failure;
	assert RAM(20136) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(20136))))  severity failure;
	assert RAM(20137) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20137))))  severity failure;
	assert RAM(20138) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(20138))))  severity failure;
	assert RAM(20139) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(20139))))  severity failure;
	assert RAM(20140) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(20140))))  severity failure;
	assert RAM(20141) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20141))))  severity failure;
	assert RAM(20142) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(20142))))  severity failure;
	assert RAM(20143) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(20143))))  severity failure;
	assert RAM(20144) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(20144))))  severity failure;
	assert RAM(20145) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20145))))  severity failure;
	assert RAM(20146) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(20146))))  severity failure;
	assert RAM(20147) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(20147))))  severity failure;
	assert RAM(20148) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(20148))))  severity failure;
	assert RAM(20149) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(20149))))  severity failure;
	assert RAM(20150) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20150))))  severity failure;
	assert RAM(20151) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(20151))))  severity failure;
	assert RAM(20152) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(20152))))  severity failure;
	assert RAM(20153) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(20153))))  severity failure;
	assert RAM(20154) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(20154))))  severity failure;
	assert RAM(20155) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(20155))))  severity failure;
	assert RAM(20156) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20156))))  severity failure;
	assert RAM(20157) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(20157))))  severity failure;
	assert RAM(20158) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(20158))))  severity failure;
	assert RAM(20159) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20159))))  severity failure;
	assert RAM(20160) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(20160))))  severity failure;
	assert RAM(20161) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(20161))))  severity failure;
	assert RAM(20162) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20162))))  severity failure;
	assert RAM(20163) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(20163))))  severity failure;
	assert RAM(20164) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20164))))  severity failure;
	assert RAM(20165) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20165))))  severity failure;
	assert RAM(20166) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(20166))))  severity failure;
	assert RAM(20167) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(20167))))  severity failure;
	assert RAM(20168) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(20168))))  severity failure;
	assert RAM(20169) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(20169))))  severity failure;
	assert RAM(20170) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20170))))  severity failure;
	assert RAM(20171) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(20171))))  severity failure;
	assert RAM(20172) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20172))))  severity failure;
	assert RAM(20173) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(20173))))  severity failure;
	assert RAM(20174) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(20174))))  severity failure;
	assert RAM(20175) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20175))))  severity failure;
	assert RAM(20176) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(20176))))  severity failure;
	assert RAM(20177) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(20177))))  severity failure;
	assert RAM(20178) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(20178))))  severity failure;
	assert RAM(20179) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(20179))))  severity failure;
	assert RAM(20180) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20180))))  severity failure;
	assert RAM(20181) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(20181))))  severity failure;
	assert RAM(20182) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(20182))))  severity failure;
	assert RAM(20183) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(20183))))  severity failure;
	assert RAM(20184) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(20184))))  severity failure;
	assert RAM(20185) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(20185))))  severity failure;
	assert RAM(20186) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(20186))))  severity failure;
	assert RAM(20187) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(20187))))  severity failure;
	assert RAM(20188) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20188))))  severity failure;
	assert RAM(20189) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20189))))  severity failure;
	assert RAM(20190) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(20190))))  severity failure;
	assert RAM(20191) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(20191))))  severity failure;
	assert RAM(20192) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(20192))))  severity failure;
	assert RAM(20193) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(20193))))  severity failure;
	assert RAM(20194) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20194))))  severity failure;
	assert RAM(20195) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20195))))  severity failure;
	assert RAM(20196) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(20196))))  severity failure;
	assert RAM(20197) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(20197))))  severity failure;
	assert RAM(20198) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20198))))  severity failure;
	assert RAM(20199) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(20199))))  severity failure;
	assert RAM(20200) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(20200))))  severity failure;
	assert RAM(20201) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(20201))))  severity failure;
	assert RAM(20202) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20202))))  severity failure;
	assert RAM(20203) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(20203))))  severity failure;
	assert RAM(20204) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(20204))))  severity failure;
	assert RAM(20205) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20205))))  severity failure;
	assert RAM(20206) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(20206))))  severity failure;
	assert RAM(20207) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(20207))))  severity failure;
	assert RAM(20208) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(20208))))  severity failure;
	assert RAM(20209) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20209))))  severity failure;
	assert RAM(20210) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(20210))))  severity failure;
	assert RAM(20211) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20211))))  severity failure;
	assert RAM(20212) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20212))))  severity failure;
	assert RAM(20213) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20213))))  severity failure;
	assert RAM(20214) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20214))))  severity failure;
	assert RAM(20215) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(20215))))  severity failure;
	assert RAM(20216) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20216))))  severity failure;
	assert RAM(20217) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(20217))))  severity failure;
	assert RAM(20218) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(20218))))  severity failure;
	assert RAM(20219) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20219))))  severity failure;
	assert RAM(20220) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(20220))))  severity failure;
	assert RAM(20221) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20221))))  severity failure;
	assert RAM(20222) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20222))))  severity failure;
	assert RAM(20223) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(20223))))  severity failure;
	assert RAM(20224) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(20224))))  severity failure;
	assert RAM(20225) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20225))))  severity failure;
	assert RAM(20226) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20226))))  severity failure;
	assert RAM(20227) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(20227))))  severity failure;
	assert RAM(20228) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(20228))))  severity failure;
	assert RAM(20229) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20229))))  severity failure;
	assert RAM(20230) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(20230))))  severity failure;
	assert RAM(20231) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20231))))  severity failure;
	assert RAM(20232) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(20232))))  severity failure;
	assert RAM(20233) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20233))))  severity failure;
	assert RAM(20234) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(20234))))  severity failure;
	assert RAM(20235) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(20235))))  severity failure;
	assert RAM(20236) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(20236))))  severity failure;
	assert RAM(20237) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20237))))  severity failure;
	assert RAM(20238) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(20238))))  severity failure;
	assert RAM(20239) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(20239))))  severity failure;
	assert RAM(20240) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(20240))))  severity failure;
	assert RAM(20241) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(20241))))  severity failure;
	assert RAM(20242) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(20242))))  severity failure;
	assert RAM(20243) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(20243))))  severity failure;
	assert RAM(20244) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(20244))))  severity failure;
	assert RAM(20245) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(20245))))  severity failure;
	assert RAM(20246) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(20246))))  severity failure;
	assert RAM(20247) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(20247))))  severity failure;
	assert RAM(20248) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(20248))))  severity failure;
	assert RAM(20249) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(20249))))  severity failure;
	assert RAM(20250) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(20250))))  severity failure;
	assert RAM(20251) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20251))))  severity failure;
	assert RAM(20252) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(20252))))  severity failure;
	assert RAM(20253) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20253))))  severity failure;
	assert RAM(20254) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(20254))))  severity failure;
	assert RAM(20255) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(20255))))  severity failure;
	assert RAM(20256) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20256))))  severity failure;
	assert RAM(20257) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(20257))))  severity failure;
	assert RAM(20258) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(20258))))  severity failure;
	assert RAM(20259) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(20259))))  severity failure;
	assert RAM(20260) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(20260))))  severity failure;
	assert RAM(20261) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20261))))  severity failure;
	assert RAM(20262) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(20262))))  severity failure;
	assert RAM(20263) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(20263))))  severity failure;
	assert RAM(20264) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20264))))  severity failure;
	assert RAM(20265) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20265))))  severity failure;
	assert RAM(20266) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20266))))  severity failure;
	assert RAM(20267) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20267))))  severity failure;
	assert RAM(20268) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(20268))))  severity failure;
	assert RAM(20269) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20269))))  severity failure;
	assert RAM(20270) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20270))))  severity failure;
	assert RAM(20271) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(20271))))  severity failure;
	assert RAM(20272) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(20272))))  severity failure;
	assert RAM(20273) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20273))))  severity failure;
	assert RAM(20274) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(20274))))  severity failure;
	assert RAM(20275) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(20275))))  severity failure;
	assert RAM(20276) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20276))))  severity failure;
	assert RAM(20277) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(20277))))  severity failure;
	assert RAM(20278) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(20278))))  severity failure;
	assert RAM(20279) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20279))))  severity failure;
	assert RAM(20280) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20280))))  severity failure;
	assert RAM(20281) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(20281))))  severity failure;
	assert RAM(20282) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20282))))  severity failure;
	assert RAM(20283) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(20283))))  severity failure;
	assert RAM(20284) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20284))))  severity failure;
	assert RAM(20285) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(20285))))  severity failure;
	assert RAM(20286) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(20286))))  severity failure;
	assert RAM(20287) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20287))))  severity failure;
	assert RAM(20288) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(20288))))  severity failure;
	assert RAM(20289) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20289))))  severity failure;
	assert RAM(20290) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(20290))))  severity failure;
	assert RAM(20291) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(20291))))  severity failure;
	assert RAM(20292) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(20292))))  severity failure;
	assert RAM(20293) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20293))))  severity failure;
	assert RAM(20294) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20294))))  severity failure;
	assert RAM(20295) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(20295))))  severity failure;
	assert RAM(20296) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(20296))))  severity failure;
	assert RAM(20297) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(20297))))  severity failure;
	assert RAM(20298) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(20298))))  severity failure;
	assert RAM(20299) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20299))))  severity failure;
	assert RAM(20300) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(20300))))  severity failure;
	assert RAM(20301) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20301))))  severity failure;
	assert RAM(20302) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(20302))))  severity failure;
	assert RAM(20303) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(20303))))  severity failure;
	assert RAM(20304) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20304))))  severity failure;
	assert RAM(20305) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20305))))  severity failure;
	assert RAM(20306) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(20306))))  severity failure;
	assert RAM(20307) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20307))))  severity failure;
	assert RAM(20308) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(20308))))  severity failure;
	assert RAM(20309) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20309))))  severity failure;
	assert RAM(20310) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(20310))))  severity failure;
	assert RAM(20311) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(20311))))  severity failure;
	assert RAM(20312) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(20312))))  severity failure;
	assert RAM(20313) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20313))))  severity failure;
	assert RAM(20314) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(20314))))  severity failure;
	assert RAM(20315) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(20315))))  severity failure;
	assert RAM(20316) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(20316))))  severity failure;
	assert RAM(20317) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(20317))))  severity failure;
	assert RAM(20318) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(20318))))  severity failure;
	assert RAM(20319) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(20319))))  severity failure;
	assert RAM(20320) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(20320))))  severity failure;
	assert RAM(20321) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(20321))))  severity failure;
	assert RAM(20322) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(20322))))  severity failure;
	assert RAM(20323) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20323))))  severity failure;
	assert RAM(20324) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20324))))  severity failure;
	assert RAM(20325) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20325))))  severity failure;
	assert RAM(20326) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(20326))))  severity failure;
	assert RAM(20327) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(20327))))  severity failure;
	assert RAM(20328) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(20328))))  severity failure;
	assert RAM(20329) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20329))))  severity failure;
	assert RAM(20330) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20330))))  severity failure;
	assert RAM(20331) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20331))))  severity failure;
	assert RAM(20332) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(20332))))  severity failure;
	assert RAM(20333) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(20333))))  severity failure;
	assert RAM(20334) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(20334))))  severity failure;
	assert RAM(20335) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(20335))))  severity failure;
	assert RAM(20336) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20336))))  severity failure;
	assert RAM(20337) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(20337))))  severity failure;
	assert RAM(20338) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(20338))))  severity failure;
	assert RAM(20339) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20339))))  severity failure;
	assert RAM(20340) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(20340))))  severity failure;
	assert RAM(20341) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(20341))))  severity failure;
	assert RAM(20342) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(20342))))  severity failure;
	assert RAM(20343) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(20343))))  severity failure;
	assert RAM(20344) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20344))))  severity failure;
	assert RAM(20345) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(20345))))  severity failure;
	assert RAM(20346) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(20346))))  severity failure;
	assert RAM(20347) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20347))))  severity failure;
	assert RAM(20348) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(20348))))  severity failure;
	assert RAM(20349) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(20349))))  severity failure;
	assert RAM(20350) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20350))))  severity failure;
	assert RAM(20351) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(20351))))  severity failure;
	assert RAM(20352) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(20352))))  severity failure;
	assert RAM(20353) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(20353))))  severity failure;
	assert RAM(20354) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20354))))  severity failure;
	assert RAM(20355) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(20355))))  severity failure;
	assert RAM(20356) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(20356))))  severity failure;
	assert RAM(20357) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(20357))))  severity failure;
	assert RAM(20358) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(20358))))  severity failure;
	assert RAM(20359) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(20359))))  severity failure;
	assert RAM(20360) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(20360))))  severity failure;
	assert RAM(20361) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(20361))))  severity failure;
	assert RAM(20362) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(20362))))  severity failure;
	assert RAM(20363) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(20363))))  severity failure;
	assert RAM(20364) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(20364))))  severity failure;
	assert RAM(20365) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(20365))))  severity failure;
	assert RAM(20366) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(20366))))  severity failure;
	assert RAM(20367) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20367))))  severity failure;
	assert RAM(20368) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20368))))  severity failure;
	assert RAM(20369) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20369))))  severity failure;
	assert RAM(20370) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(20370))))  severity failure;
	assert RAM(20371) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(20371))))  severity failure;
	assert RAM(20372) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20372))))  severity failure;
	assert RAM(20373) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(20373))))  severity failure;
	assert RAM(20374) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20374))))  severity failure;
	assert RAM(20375) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(20375))))  severity failure;
	assert RAM(20376) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(20376))))  severity failure;
	assert RAM(20377) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(20377))))  severity failure;
	assert RAM(20378) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(20378))))  severity failure;
	assert RAM(20379) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(20379))))  severity failure;
	assert RAM(20380) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(20380))))  severity failure;
	assert RAM(20381) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(20381))))  severity failure;
	assert RAM(20382) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20382))))  severity failure;
	assert RAM(20383) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20383))))  severity failure;
	assert RAM(20384) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20384))))  severity failure;
	assert RAM(20385) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20385))))  severity failure;
	assert RAM(20386) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(20386))))  severity failure;
	assert RAM(20387) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20387))))  severity failure;
	assert RAM(20388) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(20388))))  severity failure;
	assert RAM(20389) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(20389))))  severity failure;
	assert RAM(20390) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(20390))))  severity failure;
	assert RAM(20391) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20391))))  severity failure;
	assert RAM(20392) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(20392))))  severity failure;
	assert RAM(20393) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(20393))))  severity failure;
	assert RAM(20394) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(20394))))  severity failure;
	assert RAM(20395) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20395))))  severity failure;
	assert RAM(20396) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(20396))))  severity failure;
	assert RAM(20397) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(20397))))  severity failure;
	assert RAM(20398) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(20398))))  severity failure;
	assert RAM(20399) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(20399))))  severity failure;
	assert RAM(20400) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(20400))))  severity failure;
	assert RAM(20401) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20401))))  severity failure;
	assert RAM(20402) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(20402))))  severity failure;
	assert RAM(20403) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(20403))))  severity failure;
	assert RAM(20404) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(20404))))  severity failure;
	assert RAM(20405) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(20405))))  severity failure;
	assert RAM(20406) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20406))))  severity failure;
	assert RAM(20407) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(20407))))  severity failure;
	assert RAM(20408) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(20408))))  severity failure;
	assert RAM(20409) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(20409))))  severity failure;
	assert RAM(20410) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(20410))))  severity failure;
	assert RAM(20411) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(20411))))  severity failure;
	assert RAM(20412) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(20412))))  severity failure;
	assert RAM(20413) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(20413))))  severity failure;
	assert RAM(20414) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20414))))  severity failure;
	assert RAM(20415) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(20415))))  severity failure;
	assert RAM(20416) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(20416))))  severity failure;
	assert RAM(20417) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(20417))))  severity failure;
	assert RAM(20418) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(20418))))  severity failure;
	assert RAM(20419) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(20419))))  severity failure;
	assert RAM(20420) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(20420))))  severity failure;
	assert RAM(20421) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20421))))  severity failure;
	assert RAM(20422) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20422))))  severity failure;
	assert RAM(20423) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(20423))))  severity failure;
	assert RAM(20424) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(20424))))  severity failure;
	assert RAM(20425) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20425))))  severity failure;
	assert RAM(20426) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(20426))))  severity failure;
	assert RAM(20427) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20427))))  severity failure;
	assert RAM(20428) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(20428))))  severity failure;
	assert RAM(20429) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(20429))))  severity failure;
	assert RAM(20430) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(20430))))  severity failure;
	assert RAM(20431) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(20431))))  severity failure;
	assert RAM(20432) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(20432))))  severity failure;
	assert RAM(20433) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(20433))))  severity failure;
	assert RAM(20434) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(20434))))  severity failure;
	assert RAM(20435) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(20435))))  severity failure;
	assert RAM(20436) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(20436))))  severity failure;
	assert RAM(20437) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(20437))))  severity failure;
	assert RAM(20438) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(20438))))  severity failure;
	assert RAM(20439) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(20439))))  severity failure;
	assert RAM(20440) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20440))))  severity failure;
	assert RAM(20441) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(20441))))  severity failure;
	assert RAM(20442) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20442))))  severity failure;
	assert RAM(20443) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(20443))))  severity failure;
	assert RAM(20444) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(20444))))  severity failure;
	assert RAM(20445) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(20445))))  severity failure;
	assert RAM(20446) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20446))))  severity failure;
	assert RAM(20447) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20447))))  severity failure;
	assert RAM(20448) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20448))))  severity failure;
	assert RAM(20449) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(20449))))  severity failure;
	assert RAM(20450) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(20450))))  severity failure;
	assert RAM(20451) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(20451))))  severity failure;
	assert RAM(20452) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(20452))))  severity failure;
	assert RAM(20453) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(20453))))  severity failure;
	assert RAM(20454) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(20454))))  severity failure;
	assert RAM(20455) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20455))))  severity failure;
	assert RAM(20456) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20456))))  severity failure;
	assert RAM(20457) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(20457))))  severity failure;
	assert RAM(20458) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20458))))  severity failure;
	assert RAM(20459) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(20459))))  severity failure;
	assert RAM(20460) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(20460))))  severity failure;
	assert RAM(20461) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(20461))))  severity failure;
	assert RAM(20462) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(20462))))  severity failure;
	assert RAM(20463) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(20463))))  severity failure;
	assert RAM(20464) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20464))))  severity failure;
	assert RAM(20465) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20465))))  severity failure;
	assert RAM(20466) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(20466))))  severity failure;
	assert RAM(20467) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20467))))  severity failure;
	assert RAM(20468) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20468))))  severity failure;
	assert RAM(20469) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20469))))  severity failure;
	assert RAM(20470) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20470))))  severity failure;
	assert RAM(20471) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(20471))))  severity failure;
	assert RAM(20472) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(20472))))  severity failure;
	assert RAM(20473) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(20473))))  severity failure;
	assert RAM(20474) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20474))))  severity failure;
	assert RAM(20475) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(20475))))  severity failure;
	assert RAM(20476) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(20476))))  severity failure;
	assert RAM(20477) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(20477))))  severity failure;
	assert RAM(20478) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(20478))))  severity failure;
	assert RAM(20479) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(20479))))  severity failure;
	assert RAM(20480) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(20480))))  severity failure;
	assert RAM(20481) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(20481))))  severity failure;
	assert RAM(20482) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20482))))  severity failure;
	assert RAM(20483) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20483))))  severity failure;
	assert RAM(20484) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20484))))  severity failure;
	assert RAM(20485) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20485))))  severity failure;
	assert RAM(20486) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(20486))))  severity failure;
	assert RAM(20487) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(20487))))  severity failure;
	assert RAM(20488) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(20488))))  severity failure;
	assert RAM(20489) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20489))))  severity failure;
	assert RAM(20490) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(20490))))  severity failure;
	assert RAM(20491) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20491))))  severity failure;
	assert RAM(20492) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(20492))))  severity failure;
	assert RAM(20493) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20493))))  severity failure;
	assert RAM(20494) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(20494))))  severity failure;
	assert RAM(20495) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(20495))))  severity failure;
	assert RAM(20496) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(20496))))  severity failure;
	assert RAM(20497) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(20497))))  severity failure;
	assert RAM(20498) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20498))))  severity failure;
	assert RAM(20499) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(20499))))  severity failure;
	assert RAM(20500) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(20500))))  severity failure;
	assert RAM(20501) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(20501))))  severity failure;
	assert RAM(20502) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(20502))))  severity failure;
	assert RAM(20503) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(20503))))  severity failure;
	assert RAM(20504) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(20504))))  severity failure;
	assert RAM(20505) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(20505))))  severity failure;
	assert RAM(20506) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(20506))))  severity failure;
	assert RAM(20507) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(20507))))  severity failure;
	assert RAM(20508) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(20508))))  severity failure;
	assert RAM(20509) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(20509))))  severity failure;
	assert RAM(20510) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20510))))  severity failure;
	assert RAM(20511) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(20511))))  severity failure;
	assert RAM(20512) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(20512))))  severity failure;
	assert RAM(20513) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(20513))))  severity failure;
	assert RAM(20514) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(20514))))  severity failure;
	assert RAM(20515) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20515))))  severity failure;
	assert RAM(20516) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20516))))  severity failure;
	assert RAM(20517) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(20517))))  severity failure;
	assert RAM(20518) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20518))))  severity failure;
	assert RAM(20519) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(20519))))  severity failure;
	assert RAM(20520) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20520))))  severity failure;
	assert RAM(20521) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(20521))))  severity failure;
	assert RAM(20522) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20522))))  severity failure;
	assert RAM(20523) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20523))))  severity failure;
	assert RAM(20524) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(20524))))  severity failure;
	assert RAM(20525) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(20525))))  severity failure;
	assert RAM(20526) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(20526))))  severity failure;
	assert RAM(20527) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(20527))))  severity failure;
	assert RAM(20528) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20528))))  severity failure;
	assert RAM(20529) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(20529))))  severity failure;
	assert RAM(20530) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20530))))  severity failure;
	assert RAM(20531) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20531))))  severity failure;
	assert RAM(20532) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(20532))))  severity failure;
	assert RAM(20533) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(20533))))  severity failure;
	assert RAM(20534) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(20534))))  severity failure;
	assert RAM(20535) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(20535))))  severity failure;
	assert RAM(20536) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(20536))))  severity failure;
	assert RAM(20537) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(20537))))  severity failure;
	assert RAM(20538) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(20538))))  severity failure;
	assert RAM(20539) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(20539))))  severity failure;
	assert RAM(20540) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(20540))))  severity failure;
	assert RAM(20541) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20541))))  severity failure;
	assert RAM(20542) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(20542))))  severity failure;
	assert RAM(20543) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(20543))))  severity failure;
	assert RAM(20544) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20544))))  severity failure;
	assert RAM(20545) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20545))))  severity failure;
	assert RAM(20546) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(20546))))  severity failure;
	assert RAM(20547) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(20547))))  severity failure;
	assert RAM(20548) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(20548))))  severity failure;
	assert RAM(20549) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(20549))))  severity failure;
	assert RAM(20550) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(20550))))  severity failure;
	assert RAM(20551) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(20551))))  severity failure;
	assert RAM(20552) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(20552))))  severity failure;
	assert RAM(20553) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(20553))))  severity failure;
	assert RAM(20554) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(20554))))  severity failure;
	assert RAM(20555) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(20555))))  severity failure;
	assert RAM(20556) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(20556))))  severity failure;
	assert RAM(20557) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(20557))))  severity failure;
	assert RAM(20558) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(20558))))  severity failure;
	assert RAM(20559) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(20559))))  severity failure;
	assert RAM(20560) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(20560))))  severity failure;
	assert RAM(20561) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(20561))))  severity failure;
	assert RAM(20562) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(20562))))  severity failure;
	assert RAM(20563) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20563))))  severity failure;
	assert RAM(20564) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(20564))))  severity failure;
	assert RAM(20565) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(20565))))  severity failure;
	assert RAM(20566) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(20566))))  severity failure;
	assert RAM(20567) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20567))))  severity failure;
	assert RAM(20568) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(20568))))  severity failure;
	assert RAM(20569) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(20569))))  severity failure;
	assert RAM(20570) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(20570))))  severity failure;
	assert RAM(20571) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(20571))))  severity failure;
	assert RAM(20572) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20572))))  severity failure;
	assert RAM(20573) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20573))))  severity failure;
	assert RAM(20574) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(20574))))  severity failure;
	assert RAM(20575) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20575))))  severity failure;
	assert RAM(20576) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(20576))))  severity failure;
	assert RAM(20577) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20577))))  severity failure;
	assert RAM(20578) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(20578))))  severity failure;
	assert RAM(20579) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(20579))))  severity failure;
	assert RAM(20580) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(20580))))  severity failure;
	assert RAM(20581) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(20581))))  severity failure;
	assert RAM(20582) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20582))))  severity failure;
	assert RAM(20583) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20583))))  severity failure;
	assert RAM(20584) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20584))))  severity failure;
	assert RAM(20585) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(20585))))  severity failure;
	assert RAM(20586) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(20586))))  severity failure;
	assert RAM(20587) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(20587))))  severity failure;
	assert RAM(20588) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(20588))))  severity failure;
	assert RAM(20589) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(20589))))  severity failure;
	assert RAM(20590) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(20590))))  severity failure;
	assert RAM(20591) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(20591))))  severity failure;
	assert RAM(20592) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(20592))))  severity failure;
	assert RAM(20593) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(20593))))  severity failure;
	assert RAM(20594) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(20594))))  severity failure;
	assert RAM(20595) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(20595))))  severity failure;
	assert RAM(20596) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(20596))))  severity failure;
	assert RAM(20597) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20597))))  severity failure;
	assert RAM(20598) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20598))))  severity failure;
	assert RAM(20599) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(20599))))  severity failure;
	assert RAM(20600) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(20600))))  severity failure;
	assert RAM(20601) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(20601))))  severity failure;
	assert RAM(20602) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(20602))))  severity failure;
	assert RAM(20603) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(20603))))  severity failure;
	assert RAM(20604) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(20604))))  severity failure;
	assert RAM(20605) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20605))))  severity failure;
	assert RAM(20606) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20606))))  severity failure;
	assert RAM(20607) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20607))))  severity failure;
	assert RAM(20608) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20608))))  severity failure;
	assert RAM(20609) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20609))))  severity failure;
	assert RAM(20610) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(20610))))  severity failure;
	assert RAM(20611) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(20611))))  severity failure;
	assert RAM(20612) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(20612))))  severity failure;
	assert RAM(20613) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(20613))))  severity failure;
	assert RAM(20614) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(20614))))  severity failure;
	assert RAM(20615) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(20615))))  severity failure;
	assert RAM(20616) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(20616))))  severity failure;
	assert RAM(20617) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(20617))))  severity failure;
	assert RAM(20618) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(20618))))  severity failure;
	assert RAM(20619) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(20619))))  severity failure;
	assert RAM(20620) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(20620))))  severity failure;
	assert RAM(20621) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(20621))))  severity failure;
	assert RAM(20622) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(20622))))  severity failure;
	assert RAM(20623) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(20623))))  severity failure;
	assert RAM(20624) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(20624))))  severity failure;
	assert RAM(20625) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(20625))))  severity failure;
	assert RAM(20626) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(20626))))  severity failure;
	assert RAM(20627) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(20627))))  severity failure;
	assert RAM(20628) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(20628))))  severity failure;
	assert RAM(20629) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(20629))))  severity failure;
	assert RAM(20630) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(20630))))  severity failure;
	assert RAM(20631) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(20631))))  severity failure;
	assert RAM(20632) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(20632))))  severity failure;
	assert RAM(20633) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(20633))))  severity failure;
	assert RAM(20634) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(20634))))  severity failure;
	assert RAM(20635) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(20635))))  severity failure;
	assert RAM(20636) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(20636))))  severity failure;
	assert RAM(20637) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20637))))  severity failure;
	assert RAM(20638) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20638))))  severity failure;
	assert RAM(20639) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(20639))))  severity failure;
	assert RAM(20640) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20640))))  severity failure;
	assert RAM(20641) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(20641))))  severity failure;
	assert RAM(20642) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(20642))))  severity failure;
	assert RAM(20643) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(20643))))  severity failure;
	assert RAM(20644) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(20644))))  severity failure;
	assert RAM(20645) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(20645))))  severity failure;
	assert RAM(20646) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(20646))))  severity failure;
	assert RAM(20647) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(20647))))  severity failure;
	assert RAM(20648) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(20648))))  severity failure;
	assert RAM(20649) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(20649))))  severity failure;
	assert RAM(20650) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(20650))))  severity failure;
	assert RAM(20651) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(20651))))  severity failure;
	assert RAM(20652) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(20652))))  severity failure;
	assert RAM(20653) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(20653))))  severity failure;
	assert RAM(20654) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20654))))  severity failure;
	assert RAM(20655) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(20655))))  severity failure;
	assert RAM(20656) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(20656))))  severity failure;
	assert RAM(20657) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(20657))))  severity failure;
	assert RAM(20658) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(20658))))  severity failure;
	assert RAM(20659) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(20659))))  severity failure;
	assert RAM(20660) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(20660))))  severity failure;
	assert RAM(20661) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(20661))))  severity failure;
	assert RAM(20662) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(20662))))  severity failure;
	assert RAM(20663) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(20663))))  severity failure;
	assert RAM(20664) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(20664))))  severity failure;
	assert RAM(20665) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(20665))))  severity failure;
	assert RAM(20666) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20666))))  severity failure;
	assert RAM(20667) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(20667))))  severity failure;
	assert RAM(20668) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(20668))))  severity failure;
	assert RAM(20669) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20669))))  severity failure;
	assert RAM(20670) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(20670))))  severity failure;
	assert RAM(20671) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(20671))))  severity failure;
	assert RAM(20672) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(20672))))  severity failure;
	assert RAM(20673) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(20673))))  severity failure;
	assert RAM(20674) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20674))))  severity failure;
	assert RAM(20675) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(20675))))  severity failure;
	assert RAM(20676) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20676))))  severity failure;
	assert RAM(20677) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(20677))))  severity failure;
	assert RAM(20678) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(20678))))  severity failure;
	assert RAM(20679) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(20679))))  severity failure;
	assert RAM(20680) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(20680))))  severity failure;
	assert RAM(20681) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(20681))))  severity failure;
	assert RAM(20682) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(20682))))  severity failure;
	assert RAM(20683) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(20683))))  severity failure;
	assert RAM(20684) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20684))))  severity failure;
	assert RAM(20685) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(20685))))  severity failure;
	assert RAM(20686) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(20686))))  severity failure;
	assert RAM(20687) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(20687))))  severity failure;
	assert RAM(20688) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(20688))))  severity failure;
	assert RAM(20689) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(20689))))  severity failure;
	assert RAM(20690) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(20690))))  severity failure;
	assert RAM(20691) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(20691))))  severity failure;
	assert RAM(20692) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(20692))))  severity failure;
	assert RAM(20693) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(20693))))  severity failure;
	assert RAM(20694) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(20694))))  severity failure;
	assert RAM(20695) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20695))))  severity failure;
	assert RAM(20696) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20696))))  severity failure;
	assert RAM(20697) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(20697))))  severity failure;
	assert RAM(20698) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(20698))))  severity failure;
	assert RAM(20699) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(20699))))  severity failure;
	assert RAM(20700) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(20700))))  severity failure;
	assert RAM(20701) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(20701))))  severity failure;
	assert RAM(20702) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(20702))))  severity failure;
	assert RAM(20703) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20703))))  severity failure;
	assert RAM(20704) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(20704))))  severity failure;
	assert RAM(20705) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(20705))))  severity failure;
	assert RAM(20706) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(20706))))  severity failure;
	assert RAM(20707) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(20707))))  severity failure;
	assert RAM(20708) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(20708))))  severity failure;
	assert RAM(20709) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(20709))))  severity failure;
	assert RAM(20710) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20710))))  severity failure;
	assert RAM(20711) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(20711))))  severity failure;
	assert RAM(20712) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(20712))))  severity failure;
	assert RAM(20713) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20713))))  severity failure;
	assert RAM(20714) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(20714))))  severity failure;
	assert RAM(20715) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20715))))  severity failure;
	assert RAM(20716) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(20716))))  severity failure;
	assert RAM(20717) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(20717))))  severity failure;
	assert RAM(20718) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(20718))))  severity failure;
	assert RAM(20719) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(20719))))  severity failure;
	assert RAM(20720) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(20720))))  severity failure;
	assert RAM(20721) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(20721))))  severity failure;
	assert RAM(20722) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(20722))))  severity failure;
	assert RAM(20723) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20723))))  severity failure;
	assert RAM(20724) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(20724))))  severity failure;
	assert RAM(20725) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(20725))))  severity failure;
	assert RAM(20726) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(20726))))  severity failure;
	assert RAM(20727) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(20727))))  severity failure;
	assert RAM(20728) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(20728))))  severity failure;
	assert RAM(20729) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20729))))  severity failure;
	assert RAM(20730) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20730))))  severity failure;
	assert RAM(20731) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(20731))))  severity failure;
	assert RAM(20732) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(20732))))  severity failure;
	assert RAM(20733) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(20733))))  severity failure;
	assert RAM(20734) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(20734))))  severity failure;
	assert RAM(20735) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(20735))))  severity failure;
	assert RAM(20736) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20736))))  severity failure;
	assert RAM(20737) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(20737))))  severity failure;
	assert RAM(20738) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(20738))))  severity failure;
	assert RAM(20739) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(20739))))  severity failure;
	assert RAM(20740) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(20740))))  severity failure;
	assert RAM(20741) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(20741))))  severity failure;
	assert RAM(20742) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20742))))  severity failure;
	assert RAM(20743) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(20743))))  severity failure;
	assert RAM(20744) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(20744))))  severity failure;
	assert RAM(20745) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(20745))))  severity failure;
	assert RAM(20746) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20746))))  severity failure;
	assert RAM(20747) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(20747))))  severity failure;
	assert RAM(20748) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(20748))))  severity failure;
	assert RAM(20749) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(20749))))  severity failure;
	assert RAM(20750) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(20750))))  severity failure;
	assert RAM(20751) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(20751))))  severity failure;
	assert RAM(20752) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(20752))))  severity failure;
	assert RAM(20753) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(20753))))  severity failure;
	assert RAM(20754) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(20754))))  severity failure;
	assert RAM(20755) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(20755))))  severity failure;
	assert RAM(20756) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(20756))))  severity failure;
	assert RAM(20757) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(20757))))  severity failure;
	assert RAM(20758) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(20758))))  severity failure;
	assert RAM(20759) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(20759))))  severity failure;
	assert RAM(20760) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(20760))))  severity failure;
	assert RAM(20761) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(20761))))  severity failure;
	assert RAM(20762) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(20762))))  severity failure;
	assert RAM(20763) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(20763))))  severity failure;
	assert RAM(20764) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(20764))))  severity failure;
	assert RAM(20765) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(20765))))  severity failure;
	assert RAM(20766) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(20766))))  severity failure;
	assert RAM(20767) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(20767))))  severity failure;
	assert RAM(20768) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20768))))  severity failure;
	assert RAM(20769) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(20769))))  severity failure;
	assert RAM(20770) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(20770))))  severity failure;
	assert RAM(20771) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(20771))))  severity failure;
	assert RAM(20772) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(20772))))  severity failure;
	assert RAM(20773) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(20773))))  severity failure;
	assert RAM(20774) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(20774))))  severity failure;
	assert RAM(20775) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(20775))))  severity failure;
	assert RAM(20776) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(20776))))  severity failure;
	assert RAM(20777) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(20777))))  severity failure;
	assert RAM(20778) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(20778))))  severity failure;
	assert RAM(20779) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20779))))  severity failure;
	assert RAM(20780) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(20780))))  severity failure;
	assert RAM(20781) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(20781))))  severity failure;
	assert RAM(20782) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(20782))))  severity failure;
	assert RAM(20783) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(20783))))  severity failure;
	assert RAM(20784) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(20784))))  severity failure;
	assert RAM(20785) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(20785))))  severity failure;
	assert RAM(20786) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(20786))))  severity failure;
	assert RAM(20787) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20787))))  severity failure;
	assert RAM(20788) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(20788))))  severity failure;
	assert RAM(20789) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(20789))))  severity failure;
	assert RAM(20790) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(20790))))  severity failure;
	assert RAM(20791) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(20791))))  severity failure;
	assert RAM(20792) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(20792))))  severity failure;
	assert RAM(20793) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(20793))))  severity failure;
	assert RAM(20794) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20794))))  severity failure;
	assert RAM(20795) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(20795))))  severity failure;
	assert RAM(20796) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(20796))))  severity failure;
	assert RAM(20797) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(20797))))  severity failure;
	assert RAM(20798) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(20798))))  severity failure;
	assert RAM(20799) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(20799))))  severity failure;
	assert RAM(20800) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(20800))))  severity failure;
	assert RAM(20801) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(20801))))  severity failure;
	assert RAM(20802) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(20802))))  severity failure;
	assert RAM(20803) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(20803))))  severity failure;
	assert RAM(20804) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(20804))))  severity failure;
	assert RAM(20805) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(20805))))  severity failure;
	assert RAM(20806) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(20806))))  severity failure;
	assert RAM(20807) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(20807))))  severity failure;
	assert RAM(20808) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(20808))))  severity failure;
	assert RAM(20809) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(20809))))  severity failure;
	assert RAM(20810) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(20810))))  severity failure;
	assert RAM(20811) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(20811))))  severity failure;
	assert RAM(20812) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20812))))  severity failure;
	assert RAM(20813) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(20813))))  severity failure;
	assert RAM(20814) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(20814))))  severity failure;
	assert RAM(20815) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(20815))))  severity failure;
	assert RAM(20816) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(20816))))  severity failure;
	assert RAM(20817) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20817))))  severity failure;
	assert RAM(20818) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20818))))  severity failure;
	assert RAM(20819) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(20819))))  severity failure;
	assert RAM(20820) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20820))))  severity failure;
	assert RAM(20821) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(20821))))  severity failure;
	assert RAM(20822) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20822))))  severity failure;
	assert RAM(20823) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20823))))  severity failure;
	assert RAM(20824) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(20824))))  severity failure;
	assert RAM(20825) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(20825))))  severity failure;
	assert RAM(20826) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20826))))  severity failure;
	assert RAM(20827) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(20827))))  severity failure;
	assert RAM(20828) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20828))))  severity failure;
	assert RAM(20829) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20829))))  severity failure;
	assert RAM(20830) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(20830))))  severity failure;
	assert RAM(20831) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(20831))))  severity failure;
	assert RAM(20832) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(20832))))  severity failure;
	assert RAM(20833) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(20833))))  severity failure;
	assert RAM(20834) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(20834))))  severity failure;
	assert RAM(20835) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(20835))))  severity failure;
	assert RAM(20836) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20836))))  severity failure;
	assert RAM(20837) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20837))))  severity failure;
	assert RAM(20838) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(20838))))  severity failure;
	assert RAM(20839) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(20839))))  severity failure;
	assert RAM(20840) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(20840))))  severity failure;
	assert RAM(20841) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20841))))  severity failure;
	assert RAM(20842) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20842))))  severity failure;
	assert RAM(20843) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20843))))  severity failure;
	assert RAM(20844) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(20844))))  severity failure;
	assert RAM(20845) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20845))))  severity failure;
	assert RAM(20846) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(20846))))  severity failure;
	assert RAM(20847) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(20847))))  severity failure;
	assert RAM(20848) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(20848))))  severity failure;
	assert RAM(20849) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20849))))  severity failure;
	assert RAM(20850) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(20850))))  severity failure;
	assert RAM(20851) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(20851))))  severity failure;
	assert RAM(20852) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(20852))))  severity failure;
	assert RAM(20853) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(20853))))  severity failure;
	assert RAM(20854) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(20854))))  severity failure;
	assert RAM(20855) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(20855))))  severity failure;
	assert RAM(20856) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(20856))))  severity failure;
	assert RAM(20857) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(20857))))  severity failure;
	assert RAM(20858) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(20858))))  severity failure;
	assert RAM(20859) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(20859))))  severity failure;
	assert RAM(20860) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(20860))))  severity failure;
	assert RAM(20861) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(20861))))  severity failure;
	assert RAM(20862) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(20862))))  severity failure;
	assert RAM(20863) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(20863))))  severity failure;
	assert RAM(20864) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(20864))))  severity failure;
	assert RAM(20865) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(20865))))  severity failure;
	assert RAM(20866) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20866))))  severity failure;
	assert RAM(20867) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(20867))))  severity failure;
	assert RAM(20868) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(20868))))  severity failure;
	assert RAM(20869) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(20869))))  severity failure;
	assert RAM(20870) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(20870))))  severity failure;
	assert RAM(20871) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20871))))  severity failure;
	assert RAM(20872) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(20872))))  severity failure;
	assert RAM(20873) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(20873))))  severity failure;
	assert RAM(20874) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20874))))  severity failure;
	assert RAM(20875) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20875))))  severity failure;
	assert RAM(20876) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(20876))))  severity failure;
	assert RAM(20877) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(20877))))  severity failure;
	assert RAM(20878) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(20878))))  severity failure;
	assert RAM(20879) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(20879))))  severity failure;
	assert RAM(20880) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20880))))  severity failure;
	assert RAM(20881) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(20881))))  severity failure;
	assert RAM(20882) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(20882))))  severity failure;
	assert RAM(20883) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(20883))))  severity failure;
	assert RAM(20884) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(20884))))  severity failure;
	assert RAM(20885) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(20885))))  severity failure;
	assert RAM(20886) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(20886))))  severity failure;
	assert RAM(20887) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(20887))))  severity failure;
	assert RAM(20888) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(20888))))  severity failure;
	assert RAM(20889) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(20889))))  severity failure;
	assert RAM(20890) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(20890))))  severity failure;
	assert RAM(20891) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(20891))))  severity failure;
	assert RAM(20892) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20892))))  severity failure;
	assert RAM(20893) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(20893))))  severity failure;
	assert RAM(20894) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(20894))))  severity failure;
	assert RAM(20895) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(20895))))  severity failure;
	assert RAM(20896) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(20896))))  severity failure;
	assert RAM(20897) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(20897))))  severity failure;
	assert RAM(20898) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(20898))))  severity failure;
	assert RAM(20899) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(20899))))  severity failure;
	assert RAM(20900) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20900))))  severity failure;
	assert RAM(20901) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(20901))))  severity failure;
	assert RAM(20902) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(20902))))  severity failure;
	assert RAM(20903) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(20903))))  severity failure;
	assert RAM(20904) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(20904))))  severity failure;
	assert RAM(20905) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(20905))))  severity failure;
	assert RAM(20906) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20906))))  severity failure;
	assert RAM(20907) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(20907))))  severity failure;
	assert RAM(20908) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(20908))))  severity failure;
	assert RAM(20909) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(20909))))  severity failure;
	assert RAM(20910) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(20910))))  severity failure;
	assert RAM(20911) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(20911))))  severity failure;
	assert RAM(20912) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(20912))))  severity failure;
	assert RAM(20913) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(20913))))  severity failure;
	assert RAM(20914) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(20914))))  severity failure;
	assert RAM(20915) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(20915))))  severity failure;
	assert RAM(20916) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(20916))))  severity failure;
	assert RAM(20917) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(20917))))  severity failure;
	assert RAM(20918) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(20918))))  severity failure;
	assert RAM(20919) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(20919))))  severity failure;
	assert RAM(20920) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(20920))))  severity failure;
	assert RAM(20921) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(20921))))  severity failure;
	assert RAM(20922) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(20922))))  severity failure;
	assert RAM(20923) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(20923))))  severity failure;
	assert RAM(20924) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20924))))  severity failure;
	assert RAM(20925) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(20925))))  severity failure;
	assert RAM(20926) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20926))))  severity failure;
	assert RAM(20927) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(20927))))  severity failure;
	assert RAM(20928) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(20928))))  severity failure;
	assert RAM(20929) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(20929))))  severity failure;
	assert RAM(20930) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(20930))))  severity failure;
	assert RAM(20931) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(20931))))  severity failure;
	assert RAM(20932) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(20932))))  severity failure;
	assert RAM(20933) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(20933))))  severity failure;
	assert RAM(20934) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(20934))))  severity failure;
	assert RAM(20935) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(20935))))  severity failure;
	assert RAM(20936) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(20936))))  severity failure;
	assert RAM(20937) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(20937))))  severity failure;
	assert RAM(20938) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(20938))))  severity failure;
	assert RAM(20939) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(20939))))  severity failure;
	assert RAM(20940) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(20940))))  severity failure;
	assert RAM(20941) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(20941))))  severity failure;
	assert RAM(20942) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(20942))))  severity failure;
	assert RAM(20943) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(20943))))  severity failure;
	assert RAM(20944) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(20944))))  severity failure;
	assert RAM(20945) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(20945))))  severity failure;
	assert RAM(20946) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20946))))  severity failure;
	assert RAM(20947) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(20947))))  severity failure;
	assert RAM(20948) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(20948))))  severity failure;
	assert RAM(20949) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(20949))))  severity failure;
	assert RAM(20950) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(20950))))  severity failure;
	assert RAM(20951) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(20951))))  severity failure;
	assert RAM(20952) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(20952))))  severity failure;
	assert RAM(20953) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(20953))))  severity failure;
	assert RAM(20954) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(20954))))  severity failure;
	assert RAM(20955) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(20955))))  severity failure;
	assert RAM(20956) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(20956))))  severity failure;
	assert RAM(20957) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(20957))))  severity failure;
	assert RAM(20958) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(20958))))  severity failure;
	assert RAM(20959) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(20959))))  severity failure;
	assert RAM(20960) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20960))))  severity failure;
	assert RAM(20961) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(20961))))  severity failure;
	assert RAM(20962) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(20962))))  severity failure;
	assert RAM(20963) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(20963))))  severity failure;
	assert RAM(20964) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(20964))))  severity failure;
	assert RAM(20965) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(20965))))  severity failure;
	assert RAM(20966) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(20966))))  severity failure;
	assert RAM(20967) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(20967))))  severity failure;
	assert RAM(20968) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(20968))))  severity failure;
	assert RAM(20969) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(20969))))  severity failure;
	assert RAM(20970) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(20970))))  severity failure;
	assert RAM(20971) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(20971))))  severity failure;
	assert RAM(20972) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(20972))))  severity failure;
	assert RAM(20973) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(20973))))  severity failure;
	assert RAM(20974) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(20974))))  severity failure;
	assert RAM(20975) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(20975))))  severity failure;
	assert RAM(20976) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(20976))))  severity failure;
	assert RAM(20977) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(20977))))  severity failure;
	assert RAM(20978) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(20978))))  severity failure;
	assert RAM(20979) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(20979))))  severity failure;
	assert RAM(20980) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(20980))))  severity failure;
	assert RAM(20981) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(20981))))  severity failure;
	assert RAM(20982) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(20982))))  severity failure;
	assert RAM(20983) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(20983))))  severity failure;
	assert RAM(20984) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(20984))))  severity failure;
	assert RAM(20985) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(20985))))  severity failure;
	assert RAM(20986) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(20986))))  severity failure;
	assert RAM(20987) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(20987))))  severity failure;
	assert RAM(20988) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(20988))))  severity failure;
	assert RAM(20989) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(20989))))  severity failure;
	assert RAM(20990) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(20990))))  severity failure;
	assert RAM(20991) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(20991))))  severity failure;
	assert RAM(20992) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(20992))))  severity failure;
	assert RAM(20993) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(20993))))  severity failure;
	assert RAM(20994) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(20994))))  severity failure;
	assert RAM(20995) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(20995))))  severity failure;
	assert RAM(20996) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(20996))))  severity failure;
	assert RAM(20997) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(20997))))  severity failure;
	assert RAM(20998) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(20998))))  severity failure;
	assert RAM(20999) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(20999))))  severity failure;
	assert RAM(21000) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21000))))  severity failure;
	assert RAM(21001) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(21001))))  severity failure;
	assert RAM(21002) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21002))))  severity failure;
	assert RAM(21003) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21003))))  severity failure;
	assert RAM(21004) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(21004))))  severity failure;
	assert RAM(21005) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(21005))))  severity failure;
	assert RAM(21006) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21006))))  severity failure;
	assert RAM(21007) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21007))))  severity failure;
	assert RAM(21008) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(21008))))  severity failure;
	assert RAM(21009) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(21009))))  severity failure;
	assert RAM(21010) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21010))))  severity failure;
	assert RAM(21011) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(21011))))  severity failure;
	assert RAM(21012) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(21012))))  severity failure;
	assert RAM(21013) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21013))))  severity failure;
	assert RAM(21014) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(21014))))  severity failure;
	assert RAM(21015) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(21015))))  severity failure;
	assert RAM(21016) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(21016))))  severity failure;
	assert RAM(21017) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(21017))))  severity failure;
	assert RAM(21018) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(21018))))  severity failure;
	assert RAM(21019) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(21019))))  severity failure;
	assert RAM(21020) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21020))))  severity failure;
	assert RAM(21021) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(21021))))  severity failure;
	assert RAM(21022) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(21022))))  severity failure;
	assert RAM(21023) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(21023))))  severity failure;
	assert RAM(21024) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21024))))  severity failure;
	assert RAM(21025) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21025))))  severity failure;
	assert RAM(21026) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(21026))))  severity failure;
	assert RAM(21027) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(21027))))  severity failure;
	assert RAM(21028) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21028))))  severity failure;
	assert RAM(21029) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(21029))))  severity failure;
	assert RAM(21030) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(21030))))  severity failure;
	assert RAM(21031) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(21031))))  severity failure;
	assert RAM(21032) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(21032))))  severity failure;
	assert RAM(21033) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(21033))))  severity failure;
	assert RAM(21034) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(21034))))  severity failure;
	assert RAM(21035) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(21035))))  severity failure;
	assert RAM(21036) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21036))))  severity failure;
	assert RAM(21037) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21037))))  severity failure;
	assert RAM(21038) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21038))))  severity failure;
	assert RAM(21039) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(21039))))  severity failure;
	assert RAM(21040) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21040))))  severity failure;
	assert RAM(21041) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21041))))  severity failure;
	assert RAM(21042) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(21042))))  severity failure;
	assert RAM(21043) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21043))))  severity failure;
	assert RAM(21044) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(21044))))  severity failure;
	assert RAM(21045) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(21045))))  severity failure;
	assert RAM(21046) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21046))))  severity failure;
	assert RAM(21047) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(21047))))  severity failure;
	assert RAM(21048) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(21048))))  severity failure;
	assert RAM(21049) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21049))))  severity failure;
	assert RAM(21050) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21050))))  severity failure;
	assert RAM(21051) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(21051))))  severity failure;
	assert RAM(21052) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(21052))))  severity failure;
	assert RAM(21053) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(21053))))  severity failure;
	assert RAM(21054) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(21054))))  severity failure;
	assert RAM(21055) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(21055))))  severity failure;
	assert RAM(21056) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(21056))))  severity failure;
	assert RAM(21057) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(21057))))  severity failure;
	assert RAM(21058) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(21058))))  severity failure;
	assert RAM(21059) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(21059))))  severity failure;
	assert RAM(21060) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(21060))))  severity failure;
	assert RAM(21061) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(21061))))  severity failure;
	assert RAM(21062) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21062))))  severity failure;
	assert RAM(21063) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(21063))))  severity failure;
	assert RAM(21064) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(21064))))  severity failure;
	assert RAM(21065) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(21065))))  severity failure;
	assert RAM(21066) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(21066))))  severity failure;
	assert RAM(21067) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(21067))))  severity failure;
	assert RAM(21068) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(21068))))  severity failure;
	assert RAM(21069) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(21069))))  severity failure;
	assert RAM(21070) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(21070))))  severity failure;
	assert RAM(21071) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(21071))))  severity failure;
	assert RAM(21072) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(21072))))  severity failure;
	assert RAM(21073) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(21073))))  severity failure;
	assert RAM(21074) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(21074))))  severity failure;
	assert RAM(21075) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(21075))))  severity failure;
	assert RAM(21076) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(21076))))  severity failure;
	assert RAM(21077) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(21077))))  severity failure;
	assert RAM(21078) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(21078))))  severity failure;
	assert RAM(21079) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(21079))))  severity failure;
	assert RAM(21080) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21080))))  severity failure;
	assert RAM(21081) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(21081))))  severity failure;
	assert RAM(21082) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(21082))))  severity failure;
	assert RAM(21083) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(21083))))  severity failure;
	assert RAM(21084) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(21084))))  severity failure;
	assert RAM(21085) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(21085))))  severity failure;
	assert RAM(21086) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(21086))))  severity failure;
	assert RAM(21087) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21087))))  severity failure;
	assert RAM(21088) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(21088))))  severity failure;
	assert RAM(21089) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(21089))))  severity failure;
	assert RAM(21090) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(21090))))  severity failure;
	assert RAM(21091) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(21091))))  severity failure;
	assert RAM(21092) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(21092))))  severity failure;
	assert RAM(21093) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(21093))))  severity failure;
	assert RAM(21094) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(21094))))  severity failure;
	assert RAM(21095) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(21095))))  severity failure;
	assert RAM(21096) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(21096))))  severity failure;
	assert RAM(21097) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(21097))))  severity failure;
	assert RAM(21098) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(21098))))  severity failure;
	assert RAM(21099) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21099))))  severity failure;
	assert RAM(21100) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(21100))))  severity failure;
	assert RAM(21101) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(21101))))  severity failure;
	assert RAM(21102) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(21102))))  severity failure;
	assert RAM(21103) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21103))))  severity failure;
	assert RAM(21104) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(21104))))  severity failure;
	assert RAM(21105) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(21105))))  severity failure;
	assert RAM(21106) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(21106))))  severity failure;
	assert RAM(21107) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21107))))  severity failure;
	assert RAM(21108) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(21108))))  severity failure;
	assert RAM(21109) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(21109))))  severity failure;
	assert RAM(21110) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(21110))))  severity failure;
	assert RAM(21111) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(21111))))  severity failure;
	assert RAM(21112) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(21112))))  severity failure;
	assert RAM(21113) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(21113))))  severity failure;
	assert RAM(21114) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(21114))))  severity failure;
	assert RAM(21115) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(21115))))  severity failure;
	assert RAM(21116) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21116))))  severity failure;
	assert RAM(21117) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(21117))))  severity failure;
	assert RAM(21118) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(21118))))  severity failure;
	assert RAM(21119) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(21119))))  severity failure;
	assert RAM(21120) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(21120))))  severity failure;
	assert RAM(21121) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(21121))))  severity failure;
	assert RAM(21122) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(21122))))  severity failure;
	assert RAM(21123) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(21123))))  severity failure;
	assert RAM(21124) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(21124))))  severity failure;
	assert RAM(21125) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(21125))))  severity failure;
	assert RAM(21126) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(21126))))  severity failure;
	assert RAM(21127) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(21127))))  severity failure;
	assert RAM(21128) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(21128))))  severity failure;
	assert RAM(21129) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(21129))))  severity failure;
	assert RAM(21130) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21130))))  severity failure;
	assert RAM(21131) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(21131))))  severity failure;
	assert RAM(21132) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21132))))  severity failure;
	assert RAM(21133) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(21133))))  severity failure;
	assert RAM(21134) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(21134))))  severity failure;
	assert RAM(21135) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(21135))))  severity failure;
	assert RAM(21136) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(21136))))  severity failure;
	assert RAM(21137) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(21137))))  severity failure;
	assert RAM(21138) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21138))))  severity failure;
	assert RAM(21139) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(21139))))  severity failure;
	assert RAM(21140) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21140))))  severity failure;
	assert RAM(21141) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(21141))))  severity failure;
	assert RAM(21142) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(21142))))  severity failure;
	assert RAM(21143) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(21143))))  severity failure;
	assert RAM(21144) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(21144))))  severity failure;
	assert RAM(21145) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(21145))))  severity failure;
	assert RAM(21146) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21146))))  severity failure;
	assert RAM(21147) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(21147))))  severity failure;
	assert RAM(21148) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(21148))))  severity failure;
	assert RAM(21149) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(21149))))  severity failure;
	assert RAM(21150) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(21150))))  severity failure;
	assert RAM(21151) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(21151))))  severity failure;
	assert RAM(21152) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(21152))))  severity failure;
	assert RAM(21153) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21153))))  severity failure;
	assert RAM(21154) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(21154))))  severity failure;
	assert RAM(21155) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(21155))))  severity failure;
	assert RAM(21156) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21156))))  severity failure;
	assert RAM(21157) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(21157))))  severity failure;
	assert RAM(21158) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(21158))))  severity failure;
	assert RAM(21159) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21159))))  severity failure;
	assert RAM(21160) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21160))))  severity failure;
	assert RAM(21161) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(21161))))  severity failure;
	assert RAM(21162) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(21162))))  severity failure;
	assert RAM(21163) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(21163))))  severity failure;
	assert RAM(21164) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21164))))  severity failure;
	assert RAM(21165) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(21165))))  severity failure;
	assert RAM(21166) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(21166))))  severity failure;
	assert RAM(21167) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(21167))))  severity failure;
	assert RAM(21168) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(21168))))  severity failure;
	assert RAM(21169) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(21169))))  severity failure;
	assert RAM(21170) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(21170))))  severity failure;
	assert RAM(21171) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(21171))))  severity failure;
	assert RAM(21172) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(21172))))  severity failure;
	assert RAM(21173) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21173))))  severity failure;
	assert RAM(21174) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(21174))))  severity failure;
	assert RAM(21175) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(21175))))  severity failure;
	assert RAM(21176) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21176))))  severity failure;
	assert RAM(21177) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(21177))))  severity failure;
	assert RAM(21178) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(21178))))  severity failure;
	assert RAM(21179) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21179))))  severity failure;
	assert RAM(21180) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(21180))))  severity failure;
	assert RAM(21181) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21181))))  severity failure;
	assert RAM(21182) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(21182))))  severity failure;
	assert RAM(21183) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(21183))))  severity failure;
	assert RAM(21184) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(21184))))  severity failure;
	assert RAM(21185) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(21185))))  severity failure;
	assert RAM(21186) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(21186))))  severity failure;
	assert RAM(21187) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(21187))))  severity failure;
	assert RAM(21188) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(21188))))  severity failure;
	assert RAM(21189) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21189))))  severity failure;
	assert RAM(21190) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(21190))))  severity failure;
	assert RAM(21191) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(21191))))  severity failure;
	assert RAM(21192) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(21192))))  severity failure;
	assert RAM(21193) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(21193))))  severity failure;
	assert RAM(21194) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(21194))))  severity failure;
	assert RAM(21195) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(21195))))  severity failure;
	assert RAM(21196) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21196))))  severity failure;
	assert RAM(21197) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(21197))))  severity failure;
	assert RAM(21198) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(21198))))  severity failure;
	assert RAM(21199) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(21199))))  severity failure;
	assert RAM(21200) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21200))))  severity failure;
	assert RAM(21201) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(21201))))  severity failure;
	assert RAM(21202) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(21202))))  severity failure;
	assert RAM(21203) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21203))))  severity failure;
	assert RAM(21204) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(21204))))  severity failure;
	assert RAM(21205) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(21205))))  severity failure;
	assert RAM(21206) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(21206))))  severity failure;
	assert RAM(21207) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(21207))))  severity failure;
	assert RAM(21208) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21208))))  severity failure;
	assert RAM(21209) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(21209))))  severity failure;
	assert RAM(21210) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(21210))))  severity failure;
	assert RAM(21211) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21211))))  severity failure;
	assert RAM(21212) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21212))))  severity failure;
	assert RAM(21213) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(21213))))  severity failure;
	assert RAM(21214) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(21214))))  severity failure;
	assert RAM(21215) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(21215))))  severity failure;
	assert RAM(21216) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21216))))  severity failure;
	assert RAM(21217) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(21217))))  severity failure;
	assert RAM(21218) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(21218))))  severity failure;
	assert RAM(21219) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(21219))))  severity failure;
	assert RAM(21220) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(21220))))  severity failure;
	assert RAM(21221) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(21221))))  severity failure;
	assert RAM(21222) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21222))))  severity failure;
	assert RAM(21223) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(21223))))  severity failure;
	assert RAM(21224) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21224))))  severity failure;
	assert RAM(21225) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21225))))  severity failure;
	assert RAM(21226) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(21226))))  severity failure;
	assert RAM(21227) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(21227))))  severity failure;
	assert RAM(21228) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(21228))))  severity failure;
	assert RAM(21229) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(21229))))  severity failure;
	assert RAM(21230) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(21230))))  severity failure;
	assert RAM(21231) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(21231))))  severity failure;
	assert RAM(21232) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(21232))))  severity failure;
	assert RAM(21233) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(21233))))  severity failure;
	assert RAM(21234) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21234))))  severity failure;
	assert RAM(21235) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21235))))  severity failure;
	assert RAM(21236) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(21236))))  severity failure;
	assert RAM(21237) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(21237))))  severity failure;
	assert RAM(21238) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(21238))))  severity failure;
	assert RAM(21239) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(21239))))  severity failure;
	assert RAM(21240) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21240))))  severity failure;
	assert RAM(21241) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(21241))))  severity failure;
	assert RAM(21242) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(21242))))  severity failure;
	assert RAM(21243) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(21243))))  severity failure;
	assert RAM(21244) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(21244))))  severity failure;
	assert RAM(21245) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(21245))))  severity failure;
	assert RAM(21246) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21246))))  severity failure;
	assert RAM(21247) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(21247))))  severity failure;
	assert RAM(21248) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(21248))))  severity failure;
	assert RAM(21249) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(21249))))  severity failure;
	assert RAM(21250) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(21250))))  severity failure;
	assert RAM(21251) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21251))))  severity failure;
	assert RAM(21252) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21252))))  severity failure;
	assert RAM(21253) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(21253))))  severity failure;
	assert RAM(21254) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(21254))))  severity failure;
	assert RAM(21255) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(21255))))  severity failure;
	assert RAM(21256) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(21256))))  severity failure;
	assert RAM(21257) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(21257))))  severity failure;
	assert RAM(21258) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(21258))))  severity failure;
	assert RAM(21259) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21259))))  severity failure;
	assert RAM(21260) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(21260))))  severity failure;
	assert RAM(21261) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(21261))))  severity failure;
	assert RAM(21262) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(21262))))  severity failure;
	assert RAM(21263) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21263))))  severity failure;
	assert RAM(21264) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(21264))))  severity failure;
	assert RAM(21265) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(21265))))  severity failure;
	assert RAM(21266) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(21266))))  severity failure;
	assert RAM(21267) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(21267))))  severity failure;
	assert RAM(21268) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21268))))  severity failure;
	assert RAM(21269) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(21269))))  severity failure;
	assert RAM(21270) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21270))))  severity failure;
	assert RAM(21271) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21271))))  severity failure;
	assert RAM(21272) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(21272))))  severity failure;
	assert RAM(21273) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21273))))  severity failure;
	assert RAM(21274) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(21274))))  severity failure;
	assert RAM(21275) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21275))))  severity failure;
	assert RAM(21276) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21276))))  severity failure;
	assert RAM(21277) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(21277))))  severity failure;
	assert RAM(21278) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(21278))))  severity failure;
	assert RAM(21279) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(21279))))  severity failure;
	assert RAM(21280) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(21280))))  severity failure;
	assert RAM(21281) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(21281))))  severity failure;
	assert RAM(21282) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21282))))  severity failure;
	assert RAM(21283) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(21283))))  severity failure;
	assert RAM(21284) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21284))))  severity failure;
	assert RAM(21285) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21285))))  severity failure;
	assert RAM(21286) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(21286))))  severity failure;
	assert RAM(21287) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21287))))  severity failure;
	assert RAM(21288) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(21288))))  severity failure;
	assert RAM(21289) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(21289))))  severity failure;
	assert RAM(21290) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(21290))))  severity failure;
	assert RAM(21291) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(21291))))  severity failure;
	assert RAM(21292) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(21292))))  severity failure;
	assert RAM(21293) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(21293))))  severity failure;
	assert RAM(21294) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(21294))))  severity failure;
	assert RAM(21295) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(21295))))  severity failure;
	assert RAM(21296) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(21296))))  severity failure;
	assert RAM(21297) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(21297))))  severity failure;
	assert RAM(21298) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(21298))))  severity failure;
	assert RAM(21299) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(21299))))  severity failure;
	assert RAM(21300) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21300))))  severity failure;
	assert RAM(21301) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(21301))))  severity failure;
	assert RAM(21302) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21302))))  severity failure;
	assert RAM(21303) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(21303))))  severity failure;
	assert RAM(21304) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(21304))))  severity failure;
	assert RAM(21305) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(21305))))  severity failure;
	assert RAM(21306) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(21306))))  severity failure;
	assert RAM(21307) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21307))))  severity failure;
	assert RAM(21308) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(21308))))  severity failure;
	assert RAM(21309) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(21309))))  severity failure;
	assert RAM(21310) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(21310))))  severity failure;
	assert RAM(21311) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21311))))  severity failure;
	assert RAM(21312) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(21312))))  severity failure;
	assert RAM(21313) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(21313))))  severity failure;
	assert RAM(21314) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(21314))))  severity failure;
	assert RAM(21315) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21315))))  severity failure;
	assert RAM(21316) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(21316))))  severity failure;
	assert RAM(21317) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(21317))))  severity failure;
	assert RAM(21318) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(21318))))  severity failure;
	assert RAM(21319) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(21319))))  severity failure;
	assert RAM(21320) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(21320))))  severity failure;
	assert RAM(21321) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(21321))))  severity failure;
	assert RAM(21322) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(21322))))  severity failure;
	assert RAM(21323) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(21323))))  severity failure;
	assert RAM(21324) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21324))))  severity failure;
	assert RAM(21325) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(21325))))  severity failure;
	assert RAM(21326) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(21326))))  severity failure;
	assert RAM(21327) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21327))))  severity failure;
	assert RAM(21328) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(21328))))  severity failure;
	assert RAM(21329) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21329))))  severity failure;
	assert RAM(21330) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(21330))))  severity failure;
	assert RAM(21331) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(21331))))  severity failure;
	assert RAM(21332) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(21332))))  severity failure;
	assert RAM(21333) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(21333))))  severity failure;
	assert RAM(21334) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21334))))  severity failure;
	assert RAM(21335) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(21335))))  severity failure;
	assert RAM(21336) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(21336))))  severity failure;
	assert RAM(21337) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(21337))))  severity failure;
	assert RAM(21338) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(21338))))  severity failure;
	assert RAM(21339) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(21339))))  severity failure;
	assert RAM(21340) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(21340))))  severity failure;
	assert RAM(21341) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(21341))))  severity failure;
	assert RAM(21342) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(21342))))  severity failure;
	assert RAM(21343) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(21343))))  severity failure;
	assert RAM(21344) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(21344))))  severity failure;
	assert RAM(21345) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21345))))  severity failure;
	assert RAM(21346) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(21346))))  severity failure;
	assert RAM(21347) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(21347))))  severity failure;
	assert RAM(21348) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(21348))))  severity failure;
	assert RAM(21349) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(21349))))  severity failure;
	assert RAM(21350) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(21350))))  severity failure;
	assert RAM(21351) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(21351))))  severity failure;
	assert RAM(21352) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(21352))))  severity failure;
	assert RAM(21353) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21353))))  severity failure;
	assert RAM(21354) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(21354))))  severity failure;
	assert RAM(21355) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21355))))  severity failure;
	assert RAM(21356) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21356))))  severity failure;
	assert RAM(21357) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21357))))  severity failure;
	assert RAM(21358) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(21358))))  severity failure;
	assert RAM(21359) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21359))))  severity failure;
	assert RAM(21360) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(21360))))  severity failure;
	assert RAM(21361) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(21361))))  severity failure;
	assert RAM(21362) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21362))))  severity failure;
	assert RAM(21363) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21363))))  severity failure;
	assert RAM(21364) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(21364))))  severity failure;
	assert RAM(21365) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(21365))))  severity failure;
	assert RAM(21366) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(21366))))  severity failure;
	assert RAM(21367) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(21367))))  severity failure;
	assert RAM(21368) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21368))))  severity failure;
	assert RAM(21369) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(21369))))  severity failure;
	assert RAM(21370) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(21370))))  severity failure;
	assert RAM(21371) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(21371))))  severity failure;
	assert RAM(21372) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21372))))  severity failure;
	assert RAM(21373) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21373))))  severity failure;
	assert RAM(21374) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(21374))))  severity failure;
	assert RAM(21375) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(21375))))  severity failure;
	assert RAM(21376) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(21376))))  severity failure;
	assert RAM(21377) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(21377))))  severity failure;
	assert RAM(21378) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(21378))))  severity failure;
	assert RAM(21379) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(21379))))  severity failure;
	assert RAM(21380) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21380))))  severity failure;
	assert RAM(21381) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(21381))))  severity failure;
	assert RAM(21382) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21382))))  severity failure;
	assert RAM(21383) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(21383))))  severity failure;
	assert RAM(21384) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(21384))))  severity failure;
	assert RAM(21385) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(21385))))  severity failure;
	assert RAM(21386) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21386))))  severity failure;
	assert RAM(21387) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(21387))))  severity failure;
	assert RAM(21388) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(21388))))  severity failure;
	assert RAM(21389) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(21389))))  severity failure;
	assert RAM(21390) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(21390))))  severity failure;
	assert RAM(21391) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(21391))))  severity failure;
	assert RAM(21392) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21392))))  severity failure;
	assert RAM(21393) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(21393))))  severity failure;
	assert RAM(21394) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(21394))))  severity failure;
	assert RAM(21395) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(21395))))  severity failure;
	assert RAM(21396) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(21396))))  severity failure;
	assert RAM(21397) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(21397))))  severity failure;
	assert RAM(21398) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(21398))))  severity failure;
	assert RAM(21399) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(21399))))  severity failure;
	assert RAM(21400) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(21400))))  severity failure;
	assert RAM(21401) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(21401))))  severity failure;
	assert RAM(21402) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(21402))))  severity failure;
	assert RAM(21403) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(21403))))  severity failure;
	assert RAM(21404) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(21404))))  severity failure;
	assert RAM(21405) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(21405))))  severity failure;
	assert RAM(21406) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21406))))  severity failure;
	assert RAM(21407) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(21407))))  severity failure;
	assert RAM(21408) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21408))))  severity failure;
	assert RAM(21409) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(21409))))  severity failure;
	assert RAM(21410) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21410))))  severity failure;
	assert RAM(21411) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(21411))))  severity failure;
	assert RAM(21412) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(21412))))  severity failure;
	assert RAM(21413) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21413))))  severity failure;
	assert RAM(21414) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(21414))))  severity failure;
	assert RAM(21415) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(21415))))  severity failure;
	assert RAM(21416) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(21416))))  severity failure;
	assert RAM(21417) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(21417))))  severity failure;
	assert RAM(21418) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21418))))  severity failure;
	assert RAM(21419) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(21419))))  severity failure;
	assert RAM(21420) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21420))))  severity failure;
	assert RAM(21421) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21421))))  severity failure;
	assert RAM(21422) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21422))))  severity failure;
	assert RAM(21423) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21423))))  severity failure;
	assert RAM(21424) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(21424))))  severity failure;
	assert RAM(21425) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(21425))))  severity failure;
	assert RAM(21426) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(21426))))  severity failure;
	assert RAM(21427) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(21427))))  severity failure;
	assert RAM(21428) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(21428))))  severity failure;
	assert RAM(21429) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(21429))))  severity failure;
	assert RAM(21430) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21430))))  severity failure;
	assert RAM(21431) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(21431))))  severity failure;
	assert RAM(21432) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(21432))))  severity failure;
	assert RAM(21433) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(21433))))  severity failure;
	assert RAM(21434) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(21434))))  severity failure;
	assert RAM(21435) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(21435))))  severity failure;
	assert RAM(21436) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21436))))  severity failure;
	assert RAM(21437) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(21437))))  severity failure;
	assert RAM(21438) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(21438))))  severity failure;
	assert RAM(21439) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(21439))))  severity failure;
	assert RAM(21440) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(21440))))  severity failure;
	assert RAM(21441) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21441))))  severity failure;
	assert RAM(21442) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(21442))))  severity failure;
	assert RAM(21443) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21443))))  severity failure;
	assert RAM(21444) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(21444))))  severity failure;
	assert RAM(21445) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(21445))))  severity failure;
	assert RAM(21446) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(21446))))  severity failure;
	assert RAM(21447) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(21447))))  severity failure;
	assert RAM(21448) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(21448))))  severity failure;
	assert RAM(21449) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21449))))  severity failure;
	assert RAM(21450) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(21450))))  severity failure;
	assert RAM(21451) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21451))))  severity failure;
	assert RAM(21452) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21452))))  severity failure;
	assert RAM(21453) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(21453))))  severity failure;
	assert RAM(21454) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(21454))))  severity failure;
	assert RAM(21455) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(21455))))  severity failure;
	assert RAM(21456) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(21456))))  severity failure;
	assert RAM(21457) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21457))))  severity failure;
	assert RAM(21458) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(21458))))  severity failure;
	assert RAM(21459) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(21459))))  severity failure;
	assert RAM(21460) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(21460))))  severity failure;
	assert RAM(21461) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21461))))  severity failure;
	assert RAM(21462) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21462))))  severity failure;
	assert RAM(21463) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(21463))))  severity failure;
	assert RAM(21464) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(21464))))  severity failure;
	assert RAM(21465) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(21465))))  severity failure;
	assert RAM(21466) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(21466))))  severity failure;
	assert RAM(21467) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(21467))))  severity failure;
	assert RAM(21468) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(21468))))  severity failure;
	assert RAM(21469) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(21469))))  severity failure;
	assert RAM(21470) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(21470))))  severity failure;
	assert RAM(21471) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(21471))))  severity failure;
	assert RAM(21472) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(21472))))  severity failure;
	assert RAM(21473) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21473))))  severity failure;
	assert RAM(21474) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21474))))  severity failure;
	assert RAM(21475) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(21475))))  severity failure;
	assert RAM(21476) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21476))))  severity failure;
	assert RAM(21477) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(21477))))  severity failure;
	assert RAM(21478) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(21478))))  severity failure;
	assert RAM(21479) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(21479))))  severity failure;
	assert RAM(21480) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21480))))  severity failure;
	assert RAM(21481) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(21481))))  severity failure;
	assert RAM(21482) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(21482))))  severity failure;
	assert RAM(21483) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(21483))))  severity failure;
	assert RAM(21484) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(21484))))  severity failure;
	assert RAM(21485) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(21485))))  severity failure;
	assert RAM(21486) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(21486))))  severity failure;
	assert RAM(21487) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21487))))  severity failure;
	assert RAM(21488) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(21488))))  severity failure;
	assert RAM(21489) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(21489))))  severity failure;
	assert RAM(21490) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21490))))  severity failure;
	assert RAM(21491) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(21491))))  severity failure;
	assert RAM(21492) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(21492))))  severity failure;
	assert RAM(21493) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(21493))))  severity failure;
	assert RAM(21494) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(21494))))  severity failure;
	assert RAM(21495) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21495))))  severity failure;
	assert RAM(21496) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(21496))))  severity failure;
	assert RAM(21497) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(21497))))  severity failure;
	assert RAM(21498) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(21498))))  severity failure;
	assert RAM(21499) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(21499))))  severity failure;
	assert RAM(21500) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(21500))))  severity failure;
	assert RAM(21501) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21501))))  severity failure;
	assert RAM(21502) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(21502))))  severity failure;
	assert RAM(21503) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(21503))))  severity failure;
	assert RAM(21504) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21504))))  severity failure;
	assert RAM(21505) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(21505))))  severity failure;
	assert RAM(21506) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(21506))))  severity failure;
	assert RAM(21507) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21507))))  severity failure;
	assert RAM(21508) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(21508))))  severity failure;
	assert RAM(21509) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(21509))))  severity failure;
	assert RAM(21510) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(21510))))  severity failure;
	assert RAM(21511) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(21511))))  severity failure;
	assert RAM(21512) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(21512))))  severity failure;
	assert RAM(21513) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(21513))))  severity failure;
	assert RAM(21514) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(21514))))  severity failure;
	assert RAM(21515) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21515))))  severity failure;
	assert RAM(21516) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(21516))))  severity failure;
	assert RAM(21517) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21517))))  severity failure;
	assert RAM(21518) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(21518))))  severity failure;
	assert RAM(21519) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21519))))  severity failure;
	assert RAM(21520) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(21520))))  severity failure;
	assert RAM(21521) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(21521))))  severity failure;
	assert RAM(21522) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(21522))))  severity failure;
	assert RAM(21523) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(21523))))  severity failure;
	assert RAM(21524) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(21524))))  severity failure;
	assert RAM(21525) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21525))))  severity failure;
	assert RAM(21526) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21526))))  severity failure;
	assert RAM(21527) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(21527))))  severity failure;
	assert RAM(21528) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(21528))))  severity failure;
	assert RAM(21529) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21529))))  severity failure;
	assert RAM(21530) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(21530))))  severity failure;
	assert RAM(21531) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(21531))))  severity failure;
	assert RAM(21532) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(21532))))  severity failure;
	assert RAM(21533) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21533))))  severity failure;
	assert RAM(21534) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21534))))  severity failure;
	assert RAM(21535) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21535))))  severity failure;
	assert RAM(21536) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(21536))))  severity failure;
	assert RAM(21537) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(21537))))  severity failure;
	assert RAM(21538) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(21538))))  severity failure;
	assert RAM(21539) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(21539))))  severity failure;
	assert RAM(21540) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(21540))))  severity failure;
	assert RAM(21541) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(21541))))  severity failure;
	assert RAM(21542) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(21542))))  severity failure;
	assert RAM(21543) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21543))))  severity failure;
	assert RAM(21544) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(21544))))  severity failure;
	assert RAM(21545) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21545))))  severity failure;
	assert RAM(21546) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(21546))))  severity failure;
	assert RAM(21547) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(21547))))  severity failure;
	assert RAM(21548) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(21548))))  severity failure;
	assert RAM(21549) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(21549))))  severity failure;
	assert RAM(21550) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(21550))))  severity failure;
	assert RAM(21551) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(21551))))  severity failure;
	assert RAM(21552) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(21552))))  severity failure;
	assert RAM(21553) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(21553))))  severity failure;
	assert RAM(21554) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(21554))))  severity failure;
	assert RAM(21555) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(21555))))  severity failure;
	assert RAM(21556) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21556))))  severity failure;
	assert RAM(21557) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(21557))))  severity failure;
	assert RAM(21558) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21558))))  severity failure;
	assert RAM(21559) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(21559))))  severity failure;
	assert RAM(21560) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(21560))))  severity failure;
	assert RAM(21561) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(21561))))  severity failure;
	assert RAM(21562) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(21562))))  severity failure;
	assert RAM(21563) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(21563))))  severity failure;
	assert RAM(21564) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(21564))))  severity failure;
	assert RAM(21565) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21565))))  severity failure;
	assert RAM(21566) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21566))))  severity failure;
	assert RAM(21567) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(21567))))  severity failure;
	assert RAM(21568) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(21568))))  severity failure;
	assert RAM(21569) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(21569))))  severity failure;
	assert RAM(21570) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(21570))))  severity failure;
	assert RAM(21571) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21571))))  severity failure;
	assert RAM(21572) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(21572))))  severity failure;
	assert RAM(21573) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(21573))))  severity failure;
	assert RAM(21574) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21574))))  severity failure;
	assert RAM(21575) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(21575))))  severity failure;
	assert RAM(21576) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(21576))))  severity failure;
	assert RAM(21577) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21577))))  severity failure;
	assert RAM(21578) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(21578))))  severity failure;
	assert RAM(21579) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(21579))))  severity failure;
	assert RAM(21580) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(21580))))  severity failure;
	assert RAM(21581) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21581))))  severity failure;
	assert RAM(21582) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21582))))  severity failure;
	assert RAM(21583) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(21583))))  severity failure;
	assert RAM(21584) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(21584))))  severity failure;
	assert RAM(21585) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(21585))))  severity failure;
	assert RAM(21586) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(21586))))  severity failure;
	assert RAM(21587) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(21587))))  severity failure;
	assert RAM(21588) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(21588))))  severity failure;
	assert RAM(21589) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(21589))))  severity failure;
	assert RAM(21590) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(21590))))  severity failure;
	assert RAM(21591) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(21591))))  severity failure;
	assert RAM(21592) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21592))))  severity failure;
	assert RAM(21593) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(21593))))  severity failure;
	assert RAM(21594) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(21594))))  severity failure;
	assert RAM(21595) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(21595))))  severity failure;
	assert RAM(21596) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(21596))))  severity failure;
	assert RAM(21597) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21597))))  severity failure;
	assert RAM(21598) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(21598))))  severity failure;
	assert RAM(21599) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(21599))))  severity failure;
	assert RAM(21600) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(21600))))  severity failure;
	assert RAM(21601) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(21601))))  severity failure;
	assert RAM(21602) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(21602))))  severity failure;
	assert RAM(21603) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(21603))))  severity failure;
	assert RAM(21604) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(21604))))  severity failure;
	assert RAM(21605) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(21605))))  severity failure;
	assert RAM(21606) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21606))))  severity failure;
	assert RAM(21607) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(21607))))  severity failure;
	assert RAM(21608) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(21608))))  severity failure;
	assert RAM(21609) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(21609))))  severity failure;
	assert RAM(21610) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(21610))))  severity failure;
	assert RAM(21611) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(21611))))  severity failure;
	assert RAM(21612) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(21612))))  severity failure;
	assert RAM(21613) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21613))))  severity failure;
	assert RAM(21614) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(21614))))  severity failure;
	assert RAM(21615) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(21615))))  severity failure;
	assert RAM(21616) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(21616))))  severity failure;
	assert RAM(21617) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(21617))))  severity failure;
	assert RAM(21618) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(21618))))  severity failure;
	assert RAM(21619) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21619))))  severity failure;
	assert RAM(21620) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(21620))))  severity failure;
	assert RAM(21621) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(21621))))  severity failure;
	assert RAM(21622) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(21622))))  severity failure;
	assert RAM(21623) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(21623))))  severity failure;
	assert RAM(21624) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(21624))))  severity failure;
	assert RAM(21625) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(21625))))  severity failure;
	assert RAM(21626) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(21626))))  severity failure;
	assert RAM(21627) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(21627))))  severity failure;
	assert RAM(21628) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(21628))))  severity failure;
	assert RAM(21629) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(21629))))  severity failure;
	assert RAM(21630) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(21630))))  severity failure;
	assert RAM(21631) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21631))))  severity failure;
	assert RAM(21632) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(21632))))  severity failure;
	assert RAM(21633) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(21633))))  severity failure;
	assert RAM(21634) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(21634))))  severity failure;
	assert RAM(21635) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21635))))  severity failure;
	assert RAM(21636) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(21636))))  severity failure;
	assert RAM(21637) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(21637))))  severity failure;
	assert RAM(21638) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21638))))  severity failure;
	assert RAM(21639) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(21639))))  severity failure;
	assert RAM(21640) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(21640))))  severity failure;
	assert RAM(21641) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(21641))))  severity failure;
	assert RAM(21642) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(21642))))  severity failure;
	assert RAM(21643) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(21643))))  severity failure;
	assert RAM(21644) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(21644))))  severity failure;
	assert RAM(21645) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(21645))))  severity failure;
	assert RAM(21646) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(21646))))  severity failure;
	assert RAM(21647) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(21647))))  severity failure;
	assert RAM(21648) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(21648))))  severity failure;
	assert RAM(21649) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(21649))))  severity failure;
	assert RAM(21650) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21650))))  severity failure;
	assert RAM(21651) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(21651))))  severity failure;
	assert RAM(21652) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(21652))))  severity failure;
	assert RAM(21653) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(21653))))  severity failure;
	assert RAM(21654) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(21654))))  severity failure;
	assert RAM(21655) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(21655))))  severity failure;
	assert RAM(21656) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(21656))))  severity failure;
	assert RAM(21657) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(21657))))  severity failure;
	assert RAM(21658) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(21658))))  severity failure;
	assert RAM(21659) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(21659))))  severity failure;
	assert RAM(21660) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(21660))))  severity failure;
	assert RAM(21661) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(21661))))  severity failure;
	assert RAM(21662) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(21662))))  severity failure;
	assert RAM(21663) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21663))))  severity failure;
	assert RAM(21664) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(21664))))  severity failure;
	assert RAM(21665) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(21665))))  severity failure;
	assert RAM(21666) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(21666))))  severity failure;
	assert RAM(21667) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21667))))  severity failure;
	assert RAM(21668) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(21668))))  severity failure;
	assert RAM(21669) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(21669))))  severity failure;
	assert RAM(21670) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(21670))))  severity failure;
	assert RAM(21671) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(21671))))  severity failure;
	assert RAM(21672) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(21672))))  severity failure;
	assert RAM(21673) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(21673))))  severity failure;
	assert RAM(21674) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21674))))  severity failure;
	assert RAM(21675) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(21675))))  severity failure;
	assert RAM(21676) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(21676))))  severity failure;
	assert RAM(21677) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(21677))))  severity failure;
	assert RAM(21678) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21678))))  severity failure;
	assert RAM(21679) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(21679))))  severity failure;
	assert RAM(21680) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(21680))))  severity failure;
	assert RAM(21681) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(21681))))  severity failure;
	assert RAM(21682) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(21682))))  severity failure;
	assert RAM(21683) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(21683))))  severity failure;
	assert RAM(21684) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(21684))))  severity failure;
	assert RAM(21685) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(21685))))  severity failure;
	assert RAM(21686) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21686))))  severity failure;
	assert RAM(21687) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(21687))))  severity failure;
	assert RAM(21688) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21688))))  severity failure;
	assert RAM(21689) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(21689))))  severity failure;
	assert RAM(21690) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(21690))))  severity failure;
	assert RAM(21691) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(21691))))  severity failure;
	assert RAM(21692) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21692))))  severity failure;
	assert RAM(21693) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(21693))))  severity failure;
	assert RAM(21694) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(21694))))  severity failure;
	assert RAM(21695) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(21695))))  severity failure;
	assert RAM(21696) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21696))))  severity failure;
	assert RAM(21697) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(21697))))  severity failure;
	assert RAM(21698) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(21698))))  severity failure;
	assert RAM(21699) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(21699))))  severity failure;
	assert RAM(21700) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21700))))  severity failure;
	assert RAM(21701) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(21701))))  severity failure;
	assert RAM(21702) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21702))))  severity failure;
	assert RAM(21703) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(21703))))  severity failure;
	assert RAM(21704) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(21704))))  severity failure;
	assert RAM(21705) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21705))))  severity failure;
	assert RAM(21706) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(21706))))  severity failure;
	assert RAM(21707) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(21707))))  severity failure;
	assert RAM(21708) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(21708))))  severity failure;
	assert RAM(21709) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(21709))))  severity failure;
	assert RAM(21710) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(21710))))  severity failure;
	assert RAM(21711) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21711))))  severity failure;
	assert RAM(21712) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(21712))))  severity failure;
	assert RAM(21713) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21713))))  severity failure;
	assert RAM(21714) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(21714))))  severity failure;
	assert RAM(21715) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(21715))))  severity failure;
	assert RAM(21716) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(21716))))  severity failure;
	assert RAM(21717) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(21717))))  severity failure;
	assert RAM(21718) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21718))))  severity failure;
	assert RAM(21719) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(21719))))  severity failure;
	assert RAM(21720) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(21720))))  severity failure;
	assert RAM(21721) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(21721))))  severity failure;
	assert RAM(21722) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(21722))))  severity failure;
	assert RAM(21723) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21723))))  severity failure;
	assert RAM(21724) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(21724))))  severity failure;
	assert RAM(21725) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(21725))))  severity failure;
	assert RAM(21726) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(21726))))  severity failure;
	assert RAM(21727) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21727))))  severity failure;
	assert RAM(21728) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(21728))))  severity failure;
	assert RAM(21729) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(21729))))  severity failure;
	assert RAM(21730) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(21730))))  severity failure;
	assert RAM(21731) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21731))))  severity failure;
	assert RAM(21732) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(21732))))  severity failure;
	assert RAM(21733) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(21733))))  severity failure;
	assert RAM(21734) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(21734))))  severity failure;
	assert RAM(21735) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21735))))  severity failure;
	assert RAM(21736) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(21736))))  severity failure;
	assert RAM(21737) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(21737))))  severity failure;
	assert RAM(21738) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21738))))  severity failure;
	assert RAM(21739) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(21739))))  severity failure;
	assert RAM(21740) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(21740))))  severity failure;
	assert RAM(21741) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(21741))))  severity failure;
	assert RAM(21742) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(21742))))  severity failure;
	assert RAM(21743) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(21743))))  severity failure;
	assert RAM(21744) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(21744))))  severity failure;
	assert RAM(21745) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(21745))))  severity failure;
	assert RAM(21746) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(21746))))  severity failure;
	assert RAM(21747) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(21747))))  severity failure;
	assert RAM(21748) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21748))))  severity failure;
	assert RAM(21749) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21749))))  severity failure;
	assert RAM(21750) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(21750))))  severity failure;
	assert RAM(21751) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(21751))))  severity failure;
	assert RAM(21752) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(21752))))  severity failure;
	assert RAM(21753) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(21753))))  severity failure;
	assert RAM(21754) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(21754))))  severity failure;
	assert RAM(21755) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(21755))))  severity failure;
	assert RAM(21756) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(21756))))  severity failure;
	assert RAM(21757) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(21757))))  severity failure;
	assert RAM(21758) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(21758))))  severity failure;
	assert RAM(21759) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(21759))))  severity failure;
	assert RAM(21760) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(21760))))  severity failure;
	assert RAM(21761) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(21761))))  severity failure;
	assert RAM(21762) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(21762))))  severity failure;
	assert RAM(21763) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21763))))  severity failure;
	assert RAM(21764) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(21764))))  severity failure;
	assert RAM(21765) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(21765))))  severity failure;
	assert RAM(21766) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(21766))))  severity failure;
	assert RAM(21767) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(21767))))  severity failure;
	assert RAM(21768) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(21768))))  severity failure;
	assert RAM(21769) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(21769))))  severity failure;
	assert RAM(21770) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(21770))))  severity failure;
	assert RAM(21771) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(21771))))  severity failure;
	assert RAM(21772) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(21772))))  severity failure;
	assert RAM(21773) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(21773))))  severity failure;
	assert RAM(21774) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(21774))))  severity failure;
	assert RAM(21775) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(21775))))  severity failure;
	assert RAM(21776) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(21776))))  severity failure;
	assert RAM(21777) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(21777))))  severity failure;
	assert RAM(21778) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(21778))))  severity failure;
	assert RAM(21779) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(21779))))  severity failure;
	assert RAM(21780) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21780))))  severity failure;
	assert RAM(21781) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(21781))))  severity failure;
	assert RAM(21782) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(21782))))  severity failure;
	assert RAM(21783) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(21783))))  severity failure;
	assert RAM(21784) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(21784))))  severity failure;
	assert RAM(21785) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(21785))))  severity failure;
	assert RAM(21786) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21786))))  severity failure;
	assert RAM(21787) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(21787))))  severity failure;
	assert RAM(21788) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(21788))))  severity failure;
	assert RAM(21789) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21789))))  severity failure;
	assert RAM(21790) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(21790))))  severity failure;
	assert RAM(21791) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(21791))))  severity failure;
	assert RAM(21792) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(21792))))  severity failure;
	assert RAM(21793) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21793))))  severity failure;
	assert RAM(21794) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(21794))))  severity failure;
	assert RAM(21795) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(21795))))  severity failure;
	assert RAM(21796) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(21796))))  severity failure;
	assert RAM(21797) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(21797))))  severity failure;
	assert RAM(21798) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(21798))))  severity failure;
	assert RAM(21799) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(21799))))  severity failure;
	assert RAM(21800) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(21800))))  severity failure;
	assert RAM(21801) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(21801))))  severity failure;
	assert RAM(21802) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(21802))))  severity failure;
	assert RAM(21803) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(21803))))  severity failure;
	assert RAM(21804) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21804))))  severity failure;
	assert RAM(21805) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(21805))))  severity failure;
	assert RAM(21806) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21806))))  severity failure;
	assert RAM(21807) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(21807))))  severity failure;
	assert RAM(21808) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(21808))))  severity failure;
	assert RAM(21809) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(21809))))  severity failure;
	assert RAM(21810) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(21810))))  severity failure;
	assert RAM(21811) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(21811))))  severity failure;
	assert RAM(21812) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(21812))))  severity failure;
	assert RAM(21813) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(21813))))  severity failure;
	assert RAM(21814) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21814))))  severity failure;
	assert RAM(21815) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(21815))))  severity failure;
	assert RAM(21816) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(21816))))  severity failure;
	assert RAM(21817) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(21817))))  severity failure;
	assert RAM(21818) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(21818))))  severity failure;
	assert RAM(21819) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(21819))))  severity failure;
	assert RAM(21820) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(21820))))  severity failure;
	assert RAM(21821) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(21821))))  severity failure;
	assert RAM(21822) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(21822))))  severity failure;
	assert RAM(21823) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(21823))))  severity failure;
	assert RAM(21824) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(21824))))  severity failure;
	assert RAM(21825) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(21825))))  severity failure;
	assert RAM(21826) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21826))))  severity failure;
	assert RAM(21827) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(21827))))  severity failure;
	assert RAM(21828) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(21828))))  severity failure;
	assert RAM(21829) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(21829))))  severity failure;
	assert RAM(21830) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(21830))))  severity failure;
	assert RAM(21831) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(21831))))  severity failure;
	assert RAM(21832) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(21832))))  severity failure;
	assert RAM(21833) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(21833))))  severity failure;
	assert RAM(21834) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(21834))))  severity failure;
	assert RAM(21835) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(21835))))  severity failure;
	assert RAM(21836) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(21836))))  severity failure;
	assert RAM(21837) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21837))))  severity failure;
	assert RAM(21838) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(21838))))  severity failure;
	assert RAM(21839) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(21839))))  severity failure;
	assert RAM(21840) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21840))))  severity failure;
	assert RAM(21841) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(21841))))  severity failure;
	assert RAM(21842) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(21842))))  severity failure;
	assert RAM(21843) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(21843))))  severity failure;
	assert RAM(21844) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(21844))))  severity failure;
	assert RAM(21845) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(21845))))  severity failure;
	assert RAM(21846) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21846))))  severity failure;
	assert RAM(21847) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(21847))))  severity failure;
	assert RAM(21848) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(21848))))  severity failure;
	assert RAM(21849) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21849))))  severity failure;
	assert RAM(21850) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(21850))))  severity failure;
	assert RAM(21851) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(21851))))  severity failure;
	assert RAM(21852) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(21852))))  severity failure;
	assert RAM(21853) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21853))))  severity failure;
	assert RAM(21854) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(21854))))  severity failure;
	assert RAM(21855) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(21855))))  severity failure;
	assert RAM(21856) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(21856))))  severity failure;
	assert RAM(21857) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(21857))))  severity failure;
	assert RAM(21858) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(21858))))  severity failure;
	assert RAM(21859) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(21859))))  severity failure;
	assert RAM(21860) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21860))))  severity failure;
	assert RAM(21861) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(21861))))  severity failure;
	assert RAM(21862) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(21862))))  severity failure;
	assert RAM(21863) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(21863))))  severity failure;
	assert RAM(21864) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(21864))))  severity failure;
	assert RAM(21865) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(21865))))  severity failure;
	assert RAM(21866) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21866))))  severity failure;
	assert RAM(21867) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(21867))))  severity failure;
	assert RAM(21868) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(21868))))  severity failure;
	assert RAM(21869) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(21869))))  severity failure;
	assert RAM(21870) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21870))))  severity failure;
	assert RAM(21871) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21871))))  severity failure;
	assert RAM(21872) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(21872))))  severity failure;
	assert RAM(21873) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(21873))))  severity failure;
	assert RAM(21874) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(21874))))  severity failure;
	assert RAM(21875) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(21875))))  severity failure;
	assert RAM(21876) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(21876))))  severity failure;
	assert RAM(21877) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(21877))))  severity failure;
	assert RAM(21878) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(21878))))  severity failure;
	assert RAM(21879) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(21879))))  severity failure;
	assert RAM(21880) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(21880))))  severity failure;
	assert RAM(21881) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(21881))))  severity failure;
	assert RAM(21882) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(21882))))  severity failure;
	assert RAM(21883) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(21883))))  severity failure;
	assert RAM(21884) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(21884))))  severity failure;
	assert RAM(21885) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21885))))  severity failure;
	assert RAM(21886) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(21886))))  severity failure;
	assert RAM(21887) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(21887))))  severity failure;
	assert RAM(21888) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(21888))))  severity failure;
	assert RAM(21889) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(21889))))  severity failure;
	assert RAM(21890) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(21890))))  severity failure;
	assert RAM(21891) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(21891))))  severity failure;
	assert RAM(21892) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(21892))))  severity failure;
	assert RAM(21893) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(21893))))  severity failure;
	assert RAM(21894) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(21894))))  severity failure;
	assert RAM(21895) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21895))))  severity failure;
	assert RAM(21896) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(21896))))  severity failure;
	assert RAM(21897) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(21897))))  severity failure;
	assert RAM(21898) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21898))))  severity failure;
	assert RAM(21899) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(21899))))  severity failure;
	assert RAM(21900) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(21900))))  severity failure;
	assert RAM(21901) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(21901))))  severity failure;
	assert RAM(21902) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(21902))))  severity failure;
	assert RAM(21903) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(21903))))  severity failure;
	assert RAM(21904) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(21904))))  severity failure;
	assert RAM(21905) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(21905))))  severity failure;
	assert RAM(21906) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(21906))))  severity failure;
	assert RAM(21907) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(21907))))  severity failure;
	assert RAM(21908) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(21908))))  severity failure;
	assert RAM(21909) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(21909))))  severity failure;
	assert RAM(21910) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(21910))))  severity failure;
	assert RAM(21911) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(21911))))  severity failure;
	assert RAM(21912) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(21912))))  severity failure;
	assert RAM(21913) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(21913))))  severity failure;
	assert RAM(21914) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21914))))  severity failure;
	assert RAM(21915) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(21915))))  severity failure;
	assert RAM(21916) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(21916))))  severity failure;
	assert RAM(21917) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(21917))))  severity failure;
	assert RAM(21918) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(21918))))  severity failure;
	assert RAM(21919) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(21919))))  severity failure;
	assert RAM(21920) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(21920))))  severity failure;
	assert RAM(21921) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(21921))))  severity failure;
	assert RAM(21922) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(21922))))  severity failure;
	assert RAM(21923) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(21923))))  severity failure;
	assert RAM(21924) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(21924))))  severity failure;
	assert RAM(21925) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21925))))  severity failure;
	assert RAM(21926) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(21926))))  severity failure;
	assert RAM(21927) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(21927))))  severity failure;
	assert RAM(21928) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(21928))))  severity failure;
	assert RAM(21929) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(21929))))  severity failure;
	assert RAM(21930) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(21930))))  severity failure;
	assert RAM(21931) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(21931))))  severity failure;
	assert RAM(21932) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(21932))))  severity failure;
	assert RAM(21933) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(21933))))  severity failure;
	assert RAM(21934) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(21934))))  severity failure;
	assert RAM(21935) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(21935))))  severity failure;
	assert RAM(21936) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(21936))))  severity failure;
	assert RAM(21937) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(21937))))  severity failure;
	assert RAM(21938) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(21938))))  severity failure;
	assert RAM(21939) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(21939))))  severity failure;
	assert RAM(21940) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(21940))))  severity failure;
	assert RAM(21941) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(21941))))  severity failure;
	assert RAM(21942) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(21942))))  severity failure;
	assert RAM(21943) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(21943))))  severity failure;
	assert RAM(21944) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(21944))))  severity failure;
	assert RAM(21945) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(21945))))  severity failure;
	assert RAM(21946) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(21946))))  severity failure;
	assert RAM(21947) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(21947))))  severity failure;
	assert RAM(21948) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(21948))))  severity failure;
	assert RAM(21949) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21949))))  severity failure;
	assert RAM(21950) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(21950))))  severity failure;
	assert RAM(21951) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(21951))))  severity failure;
	assert RAM(21952) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(21952))))  severity failure;
	assert RAM(21953) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(21953))))  severity failure;
	assert RAM(21954) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(21954))))  severity failure;
	assert RAM(21955) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(21955))))  severity failure;
	assert RAM(21956) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(21956))))  severity failure;
	assert RAM(21957) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(21957))))  severity failure;
	assert RAM(21958) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(21958))))  severity failure;
	assert RAM(21959) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(21959))))  severity failure;
	assert RAM(21960) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(21960))))  severity failure;
	assert RAM(21961) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(21961))))  severity failure;
	assert RAM(21962) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(21962))))  severity failure;
	assert RAM(21963) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(21963))))  severity failure;
	assert RAM(21964) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(21964))))  severity failure;
	assert RAM(21965) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(21965))))  severity failure;
	assert RAM(21966) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21966))))  severity failure;
	assert RAM(21967) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(21967))))  severity failure;
	assert RAM(21968) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(21968))))  severity failure;
	assert RAM(21969) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(21969))))  severity failure;
	assert RAM(21970) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(21970))))  severity failure;
	assert RAM(21971) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(21971))))  severity failure;
	assert RAM(21972) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21972))))  severity failure;
	assert RAM(21973) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(21973))))  severity failure;
	assert RAM(21974) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(21974))))  severity failure;
	assert RAM(21975) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(21975))))  severity failure;
	assert RAM(21976) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(21976))))  severity failure;
	assert RAM(21977) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(21977))))  severity failure;
	assert RAM(21978) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(21978))))  severity failure;
	assert RAM(21979) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(21979))))  severity failure;
	assert RAM(21980) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(21980))))  severity failure;
	assert RAM(21981) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(21981))))  severity failure;
	assert RAM(21982) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(21982))))  severity failure;
	assert RAM(21983) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(21983))))  severity failure;
	assert RAM(21984) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(21984))))  severity failure;
	assert RAM(21985) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(21985))))  severity failure;
	assert RAM(21986) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(21986))))  severity failure;
	assert RAM(21987) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(21987))))  severity failure;
	assert RAM(21988) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(21988))))  severity failure;
	assert RAM(21989) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(21989))))  severity failure;
	assert RAM(21990) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(21990))))  severity failure;
	assert RAM(21991) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(21991))))  severity failure;
	assert RAM(21992) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(21992))))  severity failure;
	assert RAM(21993) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(21993))))  severity failure;
	assert RAM(21994) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(21994))))  severity failure;
	assert RAM(21995) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(21995))))  severity failure;
	assert RAM(21996) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(21996))))  severity failure;
	assert RAM(21997) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(21997))))  severity failure;
	assert RAM(21998) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(21998))))  severity failure;
	assert RAM(21999) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(21999))))  severity failure;
	assert RAM(22000) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(22000))))  severity failure;
	assert RAM(22001) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(22001))))  severity failure;
	assert RAM(22002) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(22002))))  severity failure;
	assert RAM(22003) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(22003))))  severity failure;
	assert RAM(22004) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22004))))  severity failure;
	assert RAM(22005) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(22005))))  severity failure;
	assert RAM(22006) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(22006))))  severity failure;
	assert RAM(22007) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22007))))  severity failure;
	assert RAM(22008) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(22008))))  severity failure;
	assert RAM(22009) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(22009))))  severity failure;
	assert RAM(22010) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(22010))))  severity failure;
	assert RAM(22011) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(22011))))  severity failure;
	assert RAM(22012) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(22012))))  severity failure;
	assert RAM(22013) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(22013))))  severity failure;
	assert RAM(22014) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(22014))))  severity failure;
	assert RAM(22015) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(22015))))  severity failure;
	assert RAM(22016) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22016))))  severity failure;
	assert RAM(22017) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(22017))))  severity failure;
	assert RAM(22018) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(22018))))  severity failure;
	assert RAM(22019) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(22019))))  severity failure;
	assert RAM(22020) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(22020))))  severity failure;
	assert RAM(22021) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22021))))  severity failure;
	assert RAM(22022) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(22022))))  severity failure;
	assert RAM(22023) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(22023))))  severity failure;
	assert RAM(22024) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22024))))  severity failure;
	assert RAM(22025) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(22025))))  severity failure;
	assert RAM(22026) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(22026))))  severity failure;
	assert RAM(22027) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(22027))))  severity failure;
	assert RAM(22028) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(22028))))  severity failure;
	assert RAM(22029) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(22029))))  severity failure;
	assert RAM(22030) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(22030))))  severity failure;
	assert RAM(22031) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(22031))))  severity failure;
	assert RAM(22032) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(22032))))  severity failure;
	assert RAM(22033) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22033))))  severity failure;
	assert RAM(22034) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22034))))  severity failure;
	assert RAM(22035) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(22035))))  severity failure;
	assert RAM(22036) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(22036))))  severity failure;
	assert RAM(22037) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(22037))))  severity failure;
	assert RAM(22038) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(22038))))  severity failure;
	assert RAM(22039) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(22039))))  severity failure;
	assert RAM(22040) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(22040))))  severity failure;
	assert RAM(22041) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(22041))))  severity failure;
	assert RAM(22042) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22042))))  severity failure;
	assert RAM(22043) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22043))))  severity failure;
	assert RAM(22044) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(22044))))  severity failure;
	assert RAM(22045) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(22045))))  severity failure;
	assert RAM(22046) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(22046))))  severity failure;
	assert RAM(22047) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(22047))))  severity failure;
	assert RAM(22048) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(22048))))  severity failure;
	assert RAM(22049) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(22049))))  severity failure;
	assert RAM(22050) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(22050))))  severity failure;
	assert RAM(22051) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22051))))  severity failure;
	assert RAM(22052) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(22052))))  severity failure;
	assert RAM(22053) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(22053))))  severity failure;
	assert RAM(22054) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(22054))))  severity failure;
	assert RAM(22055) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(22055))))  severity failure;
	assert RAM(22056) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(22056))))  severity failure;
	assert RAM(22057) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(22057))))  severity failure;
	assert RAM(22058) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(22058))))  severity failure;
	assert RAM(22059) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22059))))  severity failure;
	assert RAM(22060) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22060))))  severity failure;
	assert RAM(22061) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(22061))))  severity failure;
	assert RAM(22062) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(22062))))  severity failure;
	assert RAM(22063) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(22063))))  severity failure;
	assert RAM(22064) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(22064))))  severity failure;
	assert RAM(22065) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22065))))  severity failure;
	assert RAM(22066) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(22066))))  severity failure;
	assert RAM(22067) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(22067))))  severity failure;
	assert RAM(22068) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(22068))))  severity failure;
	assert RAM(22069) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(22069))))  severity failure;
	assert RAM(22070) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22070))))  severity failure;
	assert RAM(22071) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(22071))))  severity failure;
	assert RAM(22072) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22072))))  severity failure;
	assert RAM(22073) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(22073))))  severity failure;
	assert RAM(22074) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(22074))))  severity failure;
	assert RAM(22075) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(22075))))  severity failure;
	assert RAM(22076) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22076))))  severity failure;
	assert RAM(22077) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22077))))  severity failure;
	assert RAM(22078) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(22078))))  severity failure;
	assert RAM(22079) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22079))))  severity failure;
	assert RAM(22080) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(22080))))  severity failure;
	assert RAM(22081) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(22081))))  severity failure;
	assert RAM(22082) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(22082))))  severity failure;
	assert RAM(22083) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(22083))))  severity failure;
	assert RAM(22084) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(22084))))  severity failure;
	assert RAM(22085) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22085))))  severity failure;
	assert RAM(22086) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22086))))  severity failure;
	assert RAM(22087) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(22087))))  severity failure;
	assert RAM(22088) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(22088))))  severity failure;
	assert RAM(22089) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(22089))))  severity failure;
	assert RAM(22090) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22090))))  severity failure;
	assert RAM(22091) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22091))))  severity failure;
	assert RAM(22092) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(22092))))  severity failure;
	assert RAM(22093) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(22093))))  severity failure;
	assert RAM(22094) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(22094))))  severity failure;
	assert RAM(22095) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(22095))))  severity failure;
	assert RAM(22096) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22096))))  severity failure;
	assert RAM(22097) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(22097))))  severity failure;
	assert RAM(22098) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(22098))))  severity failure;
	assert RAM(22099) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22099))))  severity failure;
	assert RAM(22100) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(22100))))  severity failure;
	assert RAM(22101) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(22101))))  severity failure;
	assert RAM(22102) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(22102))))  severity failure;
	assert RAM(22103) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22103))))  severity failure;
	assert RAM(22104) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22104))))  severity failure;
	assert RAM(22105) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(22105))))  severity failure;
	assert RAM(22106) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(22106))))  severity failure;
	assert RAM(22107) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(22107))))  severity failure;
	assert RAM(22108) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(22108))))  severity failure;
	assert RAM(22109) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(22109))))  severity failure;
	assert RAM(22110) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(22110))))  severity failure;
	assert RAM(22111) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(22111))))  severity failure;
	assert RAM(22112) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(22112))))  severity failure;
	assert RAM(22113) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(22113))))  severity failure;
	assert RAM(22114) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22114))))  severity failure;
	assert RAM(22115) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(22115))))  severity failure;
	assert RAM(22116) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(22116))))  severity failure;
	assert RAM(22117) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(22117))))  severity failure;
	assert RAM(22118) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22118))))  severity failure;
	assert RAM(22119) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22119))))  severity failure;
	assert RAM(22120) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(22120))))  severity failure;
	assert RAM(22121) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(22121))))  severity failure;
	assert RAM(22122) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22122))))  severity failure;
	assert RAM(22123) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22123))))  severity failure;
	assert RAM(22124) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22124))))  severity failure;
	assert RAM(22125) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(22125))))  severity failure;
	assert RAM(22126) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22126))))  severity failure;
	assert RAM(22127) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(22127))))  severity failure;
	assert RAM(22128) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22128))))  severity failure;
	assert RAM(22129) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(22129))))  severity failure;
	assert RAM(22130) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(22130))))  severity failure;
	assert RAM(22131) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(22131))))  severity failure;
	assert RAM(22132) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(22132))))  severity failure;
	assert RAM(22133) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22133))))  severity failure;
	assert RAM(22134) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(22134))))  severity failure;
	assert RAM(22135) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22135))))  severity failure;
	assert RAM(22136) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(22136))))  severity failure;
	assert RAM(22137) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(22137))))  severity failure;
	assert RAM(22138) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22138))))  severity failure;
	assert RAM(22139) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(22139))))  severity failure;
	assert RAM(22140) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22140))))  severity failure;
	assert RAM(22141) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(22141))))  severity failure;
	assert RAM(22142) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22142))))  severity failure;
	assert RAM(22143) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(22143))))  severity failure;
	assert RAM(22144) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(22144))))  severity failure;
	assert RAM(22145) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22145))))  severity failure;
	assert RAM(22146) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(22146))))  severity failure;
	assert RAM(22147) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(22147))))  severity failure;
	assert RAM(22148) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22148))))  severity failure;
	assert RAM(22149) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(22149))))  severity failure;
	assert RAM(22150) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(22150))))  severity failure;
	assert RAM(22151) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(22151))))  severity failure;
	assert RAM(22152) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(22152))))  severity failure;
	assert RAM(22153) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(22153))))  severity failure;
	assert RAM(22154) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(22154))))  severity failure;
	assert RAM(22155) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(22155))))  severity failure;
	assert RAM(22156) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(22156))))  severity failure;
	assert RAM(22157) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(22157))))  severity failure;
	assert RAM(22158) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(22158))))  severity failure;
	assert RAM(22159) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(22159))))  severity failure;
	assert RAM(22160) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(22160))))  severity failure;
	assert RAM(22161) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(22161))))  severity failure;
	assert RAM(22162) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(22162))))  severity failure;
	assert RAM(22163) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(22163))))  severity failure;
	assert RAM(22164) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22164))))  severity failure;
	assert RAM(22165) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(22165))))  severity failure;
	assert RAM(22166) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(22166))))  severity failure;
	assert RAM(22167) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(22167))))  severity failure;
	assert RAM(22168) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22168))))  severity failure;
	assert RAM(22169) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(22169))))  severity failure;
	assert RAM(22170) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22170))))  severity failure;
	assert RAM(22171) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(22171))))  severity failure;
	assert RAM(22172) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(22172))))  severity failure;
	assert RAM(22173) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(22173))))  severity failure;
	assert RAM(22174) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22174))))  severity failure;
	assert RAM(22175) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(22175))))  severity failure;
	assert RAM(22176) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(22176))))  severity failure;
	assert RAM(22177) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(22177))))  severity failure;
	assert RAM(22178) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(22178))))  severity failure;
	assert RAM(22179) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(22179))))  severity failure;
	assert RAM(22180) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(22180))))  severity failure;
	assert RAM(22181) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22181))))  severity failure;
	assert RAM(22182) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(22182))))  severity failure;
	assert RAM(22183) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(22183))))  severity failure;
	assert RAM(22184) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(22184))))  severity failure;
	assert RAM(22185) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22185))))  severity failure;
	assert RAM(22186) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(22186))))  severity failure;
	assert RAM(22187) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(22187))))  severity failure;
	assert RAM(22188) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22188))))  severity failure;
	assert RAM(22189) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(22189))))  severity failure;
	assert RAM(22190) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22190))))  severity failure;
	assert RAM(22191) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22191))))  severity failure;
	assert RAM(22192) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(22192))))  severity failure;
	assert RAM(22193) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(22193))))  severity failure;
	assert RAM(22194) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(22194))))  severity failure;
	assert RAM(22195) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(22195))))  severity failure;
	assert RAM(22196) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22196))))  severity failure;
	assert RAM(22197) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(22197))))  severity failure;
	assert RAM(22198) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(22198))))  severity failure;
	assert RAM(22199) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22199))))  severity failure;
	assert RAM(22200) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(22200))))  severity failure;
	assert RAM(22201) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22201))))  severity failure;
	assert RAM(22202) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(22202))))  severity failure;
	assert RAM(22203) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(22203))))  severity failure;
	assert RAM(22204) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(22204))))  severity failure;
	assert RAM(22205) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(22205))))  severity failure;
	assert RAM(22206) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(22206))))  severity failure;
	assert RAM(22207) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22207))))  severity failure;
	assert RAM(22208) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(22208))))  severity failure;
	assert RAM(22209) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(22209))))  severity failure;
	assert RAM(22210) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22210))))  severity failure;
	assert RAM(22211) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22211))))  severity failure;
	assert RAM(22212) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22212))))  severity failure;
	assert RAM(22213) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(22213))))  severity failure;
	assert RAM(22214) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(22214))))  severity failure;
	assert RAM(22215) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(22215))))  severity failure;
	assert RAM(22216) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(22216))))  severity failure;
	assert RAM(22217) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(22217))))  severity failure;
	assert RAM(22218) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(22218))))  severity failure;
	assert RAM(22219) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(22219))))  severity failure;
	assert RAM(22220) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(22220))))  severity failure;
	assert RAM(22221) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(22221))))  severity failure;
	assert RAM(22222) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(22222))))  severity failure;
	assert RAM(22223) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(22223))))  severity failure;
	assert RAM(22224) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22224))))  severity failure;
	assert RAM(22225) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(22225))))  severity failure;
	assert RAM(22226) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(22226))))  severity failure;
	assert RAM(22227) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(22227))))  severity failure;
	assert RAM(22228) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(22228))))  severity failure;
	assert RAM(22229) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22229))))  severity failure;
	assert RAM(22230) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22230))))  severity failure;
	assert RAM(22231) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(22231))))  severity failure;
	assert RAM(22232) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22232))))  severity failure;
	assert RAM(22233) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(22233))))  severity failure;
	assert RAM(22234) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22234))))  severity failure;
	assert RAM(22235) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(22235))))  severity failure;
	assert RAM(22236) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(22236))))  severity failure;
	assert RAM(22237) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22237))))  severity failure;
	assert RAM(22238) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(22238))))  severity failure;
	assert RAM(22239) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(22239))))  severity failure;
	assert RAM(22240) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(22240))))  severity failure;
	assert RAM(22241) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(22241))))  severity failure;
	assert RAM(22242) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22242))))  severity failure;
	assert RAM(22243) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22243))))  severity failure;
	assert RAM(22244) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(22244))))  severity failure;
	assert RAM(22245) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(22245))))  severity failure;
	assert RAM(22246) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(22246))))  severity failure;
	assert RAM(22247) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(22247))))  severity failure;
	assert RAM(22248) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22248))))  severity failure;
	assert RAM(22249) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(22249))))  severity failure;
	assert RAM(22250) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(22250))))  severity failure;
	assert RAM(22251) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(22251))))  severity failure;
	assert RAM(22252) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22252))))  severity failure;
	assert RAM(22253) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(22253))))  severity failure;
	assert RAM(22254) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(22254))))  severity failure;
	assert RAM(22255) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(22255))))  severity failure;
	assert RAM(22256) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(22256))))  severity failure;
	assert RAM(22257) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(22257))))  severity failure;
	assert RAM(22258) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(22258))))  severity failure;
	assert RAM(22259) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(22259))))  severity failure;
	assert RAM(22260) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(22260))))  severity failure;
	assert RAM(22261) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22261))))  severity failure;
	assert RAM(22262) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(22262))))  severity failure;
	assert RAM(22263) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(22263))))  severity failure;
	assert RAM(22264) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(22264))))  severity failure;
	assert RAM(22265) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(22265))))  severity failure;
	assert RAM(22266) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22266))))  severity failure;
	assert RAM(22267) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22267))))  severity failure;
	assert RAM(22268) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(22268))))  severity failure;
	assert RAM(22269) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22269))))  severity failure;
	assert RAM(22270) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(22270))))  severity failure;
	assert RAM(22271) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(22271))))  severity failure;
	assert RAM(22272) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(22272))))  severity failure;
	assert RAM(22273) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22273))))  severity failure;
	assert RAM(22274) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(22274))))  severity failure;
	assert RAM(22275) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(22275))))  severity failure;
	assert RAM(22276) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22276))))  severity failure;
	assert RAM(22277) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22277))))  severity failure;
	assert RAM(22278) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(22278))))  severity failure;
	assert RAM(22279) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22279))))  severity failure;
	assert RAM(22280) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22280))))  severity failure;
	assert RAM(22281) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(22281))))  severity failure;
	assert RAM(22282) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(22282))))  severity failure;
	assert RAM(22283) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(22283))))  severity failure;
	assert RAM(22284) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22284))))  severity failure;
	assert RAM(22285) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(22285))))  severity failure;
	assert RAM(22286) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(22286))))  severity failure;
	assert RAM(22287) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(22287))))  severity failure;
	assert RAM(22288) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22288))))  severity failure;
	assert RAM(22289) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(22289))))  severity failure;
	assert RAM(22290) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(22290))))  severity failure;
	assert RAM(22291) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22291))))  severity failure;
	assert RAM(22292) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(22292))))  severity failure;
	assert RAM(22293) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22293))))  severity failure;
	assert RAM(22294) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22294))))  severity failure;
	assert RAM(22295) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(22295))))  severity failure;
	assert RAM(22296) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(22296))))  severity failure;
	assert RAM(22297) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(22297))))  severity failure;
	assert RAM(22298) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(22298))))  severity failure;
	assert RAM(22299) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(22299))))  severity failure;
	assert RAM(22300) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(22300))))  severity failure;
	assert RAM(22301) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22301))))  severity failure;
	assert RAM(22302) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(22302))))  severity failure;
	assert RAM(22303) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(22303))))  severity failure;
	assert RAM(22304) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(22304))))  severity failure;
	assert RAM(22305) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(22305))))  severity failure;
	assert RAM(22306) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(22306))))  severity failure;
	assert RAM(22307) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(22307))))  severity failure;
	assert RAM(22308) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22308))))  severity failure;
	assert RAM(22309) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(22309))))  severity failure;
	assert RAM(22310) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(22310))))  severity failure;
	assert RAM(22311) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(22311))))  severity failure;
	assert RAM(22312) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(22312))))  severity failure;
	assert RAM(22313) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(22313))))  severity failure;
	assert RAM(22314) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(22314))))  severity failure;
	assert RAM(22315) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22315))))  severity failure;
	assert RAM(22316) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(22316))))  severity failure;
	assert RAM(22317) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(22317))))  severity failure;
	assert RAM(22318) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(22318))))  severity failure;
	assert RAM(22319) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(22319))))  severity failure;
	assert RAM(22320) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22320))))  severity failure;
	assert RAM(22321) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22321))))  severity failure;
	assert RAM(22322) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22322))))  severity failure;
	assert RAM(22323) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(22323))))  severity failure;
	assert RAM(22324) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(22324))))  severity failure;
	assert RAM(22325) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22325))))  severity failure;
	assert RAM(22326) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22326))))  severity failure;
	assert RAM(22327) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(22327))))  severity failure;
	assert RAM(22328) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(22328))))  severity failure;
	assert RAM(22329) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22329))))  severity failure;
	assert RAM(22330) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22330))))  severity failure;
	assert RAM(22331) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(22331))))  severity failure;
	assert RAM(22332) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(22332))))  severity failure;
	assert RAM(22333) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(22333))))  severity failure;
	assert RAM(22334) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(22334))))  severity failure;
	assert RAM(22335) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(22335))))  severity failure;
	assert RAM(22336) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(22336))))  severity failure;
	assert RAM(22337) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(22337))))  severity failure;
	assert RAM(22338) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(22338))))  severity failure;
	assert RAM(22339) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(22339))))  severity failure;
	assert RAM(22340) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(22340))))  severity failure;
	assert RAM(22341) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(22341))))  severity failure;
	assert RAM(22342) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(22342))))  severity failure;
	assert RAM(22343) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(22343))))  severity failure;
	assert RAM(22344) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(22344))))  severity failure;
	assert RAM(22345) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(22345))))  severity failure;
	assert RAM(22346) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22346))))  severity failure;
	assert RAM(22347) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22347))))  severity failure;
	assert RAM(22348) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22348))))  severity failure;
	assert RAM(22349) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(22349))))  severity failure;
	assert RAM(22350) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(22350))))  severity failure;
	assert RAM(22351) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(22351))))  severity failure;
	assert RAM(22352) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(22352))))  severity failure;
	assert RAM(22353) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(22353))))  severity failure;
	assert RAM(22354) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(22354))))  severity failure;
	assert RAM(22355) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(22355))))  severity failure;
	assert RAM(22356) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(22356))))  severity failure;
	assert RAM(22357) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(22357))))  severity failure;
	assert RAM(22358) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(22358))))  severity failure;
	assert RAM(22359) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(22359))))  severity failure;
	assert RAM(22360) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(22360))))  severity failure;
	assert RAM(22361) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(22361))))  severity failure;
	assert RAM(22362) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22362))))  severity failure;
	assert RAM(22363) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22363))))  severity failure;
	assert RAM(22364) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22364))))  severity failure;
	assert RAM(22365) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(22365))))  severity failure;
	assert RAM(22366) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(22366))))  severity failure;
	assert RAM(22367) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(22367))))  severity failure;
	assert RAM(22368) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(22368))))  severity failure;
	assert RAM(22369) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(22369))))  severity failure;
	assert RAM(22370) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(22370))))  severity failure;
	assert RAM(22371) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(22371))))  severity failure;
	assert RAM(22372) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22372))))  severity failure;
	assert RAM(22373) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22373))))  severity failure;
	assert RAM(22374) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(22374))))  severity failure;
	assert RAM(22375) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(22375))))  severity failure;
	assert RAM(22376) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(22376))))  severity failure;
	assert RAM(22377) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(22377))))  severity failure;
	assert RAM(22378) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(22378))))  severity failure;
	assert RAM(22379) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(22379))))  severity failure;
	assert RAM(22380) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(22380))))  severity failure;
	assert RAM(22381) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(22381))))  severity failure;
	assert RAM(22382) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(22382))))  severity failure;
	assert RAM(22383) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22383))))  severity failure;
	assert RAM(22384) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(22384))))  severity failure;
	assert RAM(22385) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(22385))))  severity failure;
	assert RAM(22386) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(22386))))  severity failure;
	assert RAM(22387) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22387))))  severity failure;
	assert RAM(22388) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(22388))))  severity failure;
	assert RAM(22389) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(22389))))  severity failure;
	assert RAM(22390) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(22390))))  severity failure;
	assert RAM(22391) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22391))))  severity failure;
	assert RAM(22392) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(22392))))  severity failure;
	assert RAM(22393) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22393))))  severity failure;
	assert RAM(22394) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(22394))))  severity failure;
	assert RAM(22395) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(22395))))  severity failure;
	assert RAM(22396) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(22396))))  severity failure;
	assert RAM(22397) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(22397))))  severity failure;
	assert RAM(22398) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(22398))))  severity failure;
	assert RAM(22399) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22399))))  severity failure;
	assert RAM(22400) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(22400))))  severity failure;
	assert RAM(22401) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(22401))))  severity failure;
	assert RAM(22402) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(22402))))  severity failure;
	assert RAM(22403) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(22403))))  severity failure;
	assert RAM(22404) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22404))))  severity failure;
	assert RAM(22405) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22405))))  severity failure;
	assert RAM(22406) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22406))))  severity failure;
	assert RAM(22407) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22407))))  severity failure;
	assert RAM(22408) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22408))))  severity failure;
	assert RAM(22409) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(22409))))  severity failure;
	assert RAM(22410) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(22410))))  severity failure;
	assert RAM(22411) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22411))))  severity failure;
	assert RAM(22412) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(22412))))  severity failure;
	assert RAM(22413) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(22413))))  severity failure;
	assert RAM(22414) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(22414))))  severity failure;
	assert RAM(22415) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22415))))  severity failure;
	assert RAM(22416) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(22416))))  severity failure;
	assert RAM(22417) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(22417))))  severity failure;
	assert RAM(22418) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(22418))))  severity failure;
	assert RAM(22419) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22419))))  severity failure;
	assert RAM(22420) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(22420))))  severity failure;
	assert RAM(22421) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(22421))))  severity failure;
	assert RAM(22422) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(22422))))  severity failure;
	assert RAM(22423) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(22423))))  severity failure;
	assert RAM(22424) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(22424))))  severity failure;
	assert RAM(22425) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(22425))))  severity failure;
	assert RAM(22426) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(22426))))  severity failure;
	assert RAM(22427) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(22427))))  severity failure;
	assert RAM(22428) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22428))))  severity failure;
	assert RAM(22429) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(22429))))  severity failure;
	assert RAM(22430) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22430))))  severity failure;
	assert RAM(22431) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(22431))))  severity failure;
	assert RAM(22432) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(22432))))  severity failure;
	assert RAM(22433) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22433))))  severity failure;
	assert RAM(22434) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(22434))))  severity failure;
	assert RAM(22435) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(22435))))  severity failure;
	assert RAM(22436) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22436))))  severity failure;
	assert RAM(22437) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(22437))))  severity failure;
	assert RAM(22438) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22438))))  severity failure;
	assert RAM(22439) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(22439))))  severity failure;
	assert RAM(22440) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(22440))))  severity failure;
	assert RAM(22441) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22441))))  severity failure;
	assert RAM(22442) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(22442))))  severity failure;
	assert RAM(22443) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(22443))))  severity failure;
	assert RAM(22444) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22444))))  severity failure;
	assert RAM(22445) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(22445))))  severity failure;
	assert RAM(22446) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22446))))  severity failure;
	assert RAM(22447) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22447))))  severity failure;
	assert RAM(22448) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(22448))))  severity failure;
	assert RAM(22449) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22449))))  severity failure;
	assert RAM(22450) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(22450))))  severity failure;
	assert RAM(22451) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(22451))))  severity failure;
	assert RAM(22452) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22452))))  severity failure;
	assert RAM(22453) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(22453))))  severity failure;
	assert RAM(22454) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(22454))))  severity failure;
	assert RAM(22455) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22455))))  severity failure;
	assert RAM(22456) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(22456))))  severity failure;
	assert RAM(22457) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(22457))))  severity failure;
	assert RAM(22458) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22458))))  severity failure;
	assert RAM(22459) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22459))))  severity failure;
	assert RAM(22460) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(22460))))  severity failure;
	assert RAM(22461) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22461))))  severity failure;
	assert RAM(22462) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(22462))))  severity failure;
	assert RAM(22463) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(22463))))  severity failure;
	assert RAM(22464) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(22464))))  severity failure;
	assert RAM(22465) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(22465))))  severity failure;
	assert RAM(22466) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(22466))))  severity failure;
	assert RAM(22467) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(22467))))  severity failure;
	assert RAM(22468) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(22468))))  severity failure;
	assert RAM(22469) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(22469))))  severity failure;
	assert RAM(22470) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(22470))))  severity failure;
	assert RAM(22471) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(22471))))  severity failure;
	assert RAM(22472) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(22472))))  severity failure;
	assert RAM(22473) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(22473))))  severity failure;
	assert RAM(22474) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(22474))))  severity failure;
	assert RAM(22475) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22475))))  severity failure;
	assert RAM(22476) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(22476))))  severity failure;
	assert RAM(22477) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(22477))))  severity failure;
	assert RAM(22478) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(22478))))  severity failure;
	assert RAM(22479) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22479))))  severity failure;
	assert RAM(22480) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22480))))  severity failure;
	assert RAM(22481) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22481))))  severity failure;
	assert RAM(22482) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(22482))))  severity failure;
	assert RAM(22483) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(22483))))  severity failure;
	assert RAM(22484) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(22484))))  severity failure;
	assert RAM(22485) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(22485))))  severity failure;
	assert RAM(22486) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22486))))  severity failure;
	assert RAM(22487) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(22487))))  severity failure;
	assert RAM(22488) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22488))))  severity failure;
	assert RAM(22489) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(22489))))  severity failure;
	assert RAM(22490) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(22490))))  severity failure;
	assert RAM(22491) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(22491))))  severity failure;
	assert RAM(22492) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(22492))))  severity failure;
	assert RAM(22493) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(22493))))  severity failure;
	assert RAM(22494) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(22494))))  severity failure;
	assert RAM(22495) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22495))))  severity failure;
	assert RAM(22496) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(22496))))  severity failure;
	assert RAM(22497) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(22497))))  severity failure;
	assert RAM(22498) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(22498))))  severity failure;
	assert RAM(22499) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(22499))))  severity failure;
	assert RAM(22500) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(22500))))  severity failure;
	assert RAM(22501) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(22501))))  severity failure;
	assert RAM(22502) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(22502))))  severity failure;
	assert RAM(22503) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(22503))))  severity failure;
	assert RAM(22504) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22504))))  severity failure;
	assert RAM(22505) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22505))))  severity failure;
	assert RAM(22506) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(22506))))  severity failure;
	assert RAM(22507) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(22507))))  severity failure;
	assert RAM(22508) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22508))))  severity failure;
	assert RAM(22509) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(22509))))  severity failure;
	assert RAM(22510) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(22510))))  severity failure;
	assert RAM(22511) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(22511))))  severity failure;
	assert RAM(22512) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22512))))  severity failure;
	assert RAM(22513) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(22513))))  severity failure;
	assert RAM(22514) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(22514))))  severity failure;
	assert RAM(22515) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(22515))))  severity failure;
	assert RAM(22516) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(22516))))  severity failure;
	assert RAM(22517) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22517))))  severity failure;
	assert RAM(22518) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(22518))))  severity failure;
	assert RAM(22519) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(22519))))  severity failure;
	assert RAM(22520) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22520))))  severity failure;
	assert RAM(22521) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(22521))))  severity failure;
	assert RAM(22522) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(22522))))  severity failure;
	assert RAM(22523) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(22523))))  severity failure;
	assert RAM(22524) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(22524))))  severity failure;
	assert RAM(22525) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(22525))))  severity failure;
	assert RAM(22526) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(22526))))  severity failure;
	assert RAM(22527) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(22527))))  severity failure;
	assert RAM(22528) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(22528))))  severity failure;
	assert RAM(22529) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(22529))))  severity failure;
	assert RAM(22530) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(22530))))  severity failure;
	assert RAM(22531) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(22531))))  severity failure;
	assert RAM(22532) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22532))))  severity failure;
	assert RAM(22533) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(22533))))  severity failure;
	assert RAM(22534) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22534))))  severity failure;
	assert RAM(22535) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(22535))))  severity failure;
	assert RAM(22536) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(22536))))  severity failure;
	assert RAM(22537) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(22537))))  severity failure;
	assert RAM(22538) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(22538))))  severity failure;
	assert RAM(22539) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22539))))  severity failure;
	assert RAM(22540) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22540))))  severity failure;
	assert RAM(22541) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(22541))))  severity failure;
	assert RAM(22542) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(22542))))  severity failure;
	assert RAM(22543) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(22543))))  severity failure;
	assert RAM(22544) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22544))))  severity failure;
	assert RAM(22545) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(22545))))  severity failure;
	assert RAM(22546) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(22546))))  severity failure;
	assert RAM(22547) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(22547))))  severity failure;
	assert RAM(22548) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(22548))))  severity failure;
	assert RAM(22549) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(22549))))  severity failure;
	assert RAM(22550) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22550))))  severity failure;
	assert RAM(22551) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22551))))  severity failure;
	assert RAM(22552) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22552))))  severity failure;
	assert RAM(22553) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22553))))  severity failure;
	assert RAM(22554) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22554))))  severity failure;
	assert RAM(22555) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22555))))  severity failure;
	assert RAM(22556) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(22556))))  severity failure;
	assert RAM(22557) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22557))))  severity failure;
	assert RAM(22558) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(22558))))  severity failure;
	assert RAM(22559) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(22559))))  severity failure;
	assert RAM(22560) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(22560))))  severity failure;
	assert RAM(22561) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(22561))))  severity failure;
	assert RAM(22562) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(22562))))  severity failure;
	assert RAM(22563) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(22563))))  severity failure;
	assert RAM(22564) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(22564))))  severity failure;
	assert RAM(22565) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(22565))))  severity failure;
	assert RAM(22566) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(22566))))  severity failure;
	assert RAM(22567) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22567))))  severity failure;
	assert RAM(22568) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(22568))))  severity failure;
	assert RAM(22569) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22569))))  severity failure;
	assert RAM(22570) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(22570))))  severity failure;
	assert RAM(22571) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(22571))))  severity failure;
	assert RAM(22572) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(22572))))  severity failure;
	assert RAM(22573) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(22573))))  severity failure;
	assert RAM(22574) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(22574))))  severity failure;
	assert RAM(22575) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22575))))  severity failure;
	assert RAM(22576) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(22576))))  severity failure;
	assert RAM(22577) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(22577))))  severity failure;
	assert RAM(22578) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(22578))))  severity failure;
	assert RAM(22579) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22579))))  severity failure;
	assert RAM(22580) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(22580))))  severity failure;
	assert RAM(22581) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(22581))))  severity failure;
	assert RAM(22582) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(22582))))  severity failure;
	assert RAM(22583) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(22583))))  severity failure;
	assert RAM(22584) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(22584))))  severity failure;
	assert RAM(22585) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22585))))  severity failure;
	assert RAM(22586) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(22586))))  severity failure;
	assert RAM(22587) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(22587))))  severity failure;
	assert RAM(22588) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22588))))  severity failure;
	assert RAM(22589) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(22589))))  severity failure;
	assert RAM(22590) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(22590))))  severity failure;
	assert RAM(22591) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22591))))  severity failure;
	assert RAM(22592) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(22592))))  severity failure;
	assert RAM(22593) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(22593))))  severity failure;
	assert RAM(22594) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(22594))))  severity failure;
	assert RAM(22595) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22595))))  severity failure;
	assert RAM(22596) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22596))))  severity failure;
	assert RAM(22597) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(22597))))  severity failure;
	assert RAM(22598) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(22598))))  severity failure;
	assert RAM(22599) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(22599))))  severity failure;
	assert RAM(22600) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(22600))))  severity failure;
	assert RAM(22601) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22601))))  severity failure;
	assert RAM(22602) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(22602))))  severity failure;
	assert RAM(22603) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22603))))  severity failure;
	assert RAM(22604) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(22604))))  severity failure;
	assert RAM(22605) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(22605))))  severity failure;
	assert RAM(22606) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(22606))))  severity failure;
	assert RAM(22607) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(22607))))  severity failure;
	assert RAM(22608) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(22608))))  severity failure;
	assert RAM(22609) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(22609))))  severity failure;
	assert RAM(22610) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(22610))))  severity failure;
	assert RAM(22611) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(22611))))  severity failure;
	assert RAM(22612) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(22612))))  severity failure;
	assert RAM(22613) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(22613))))  severity failure;
	assert RAM(22614) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(22614))))  severity failure;
	assert RAM(22615) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(22615))))  severity failure;
	assert RAM(22616) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(22616))))  severity failure;
	assert RAM(22617) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(22617))))  severity failure;
	assert RAM(22618) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(22618))))  severity failure;
	assert RAM(22619) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(22619))))  severity failure;
	assert RAM(22620) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22620))))  severity failure;
	assert RAM(22621) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22621))))  severity failure;
	assert RAM(22622) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22622))))  severity failure;
	assert RAM(22623) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22623))))  severity failure;
	assert RAM(22624) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(22624))))  severity failure;
	assert RAM(22625) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(22625))))  severity failure;
	assert RAM(22626) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(22626))))  severity failure;
	assert RAM(22627) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(22627))))  severity failure;
	assert RAM(22628) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22628))))  severity failure;
	assert RAM(22629) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(22629))))  severity failure;
	assert RAM(22630) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(22630))))  severity failure;
	assert RAM(22631) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(22631))))  severity failure;
	assert RAM(22632) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22632))))  severity failure;
	assert RAM(22633) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(22633))))  severity failure;
	assert RAM(22634) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(22634))))  severity failure;
	assert RAM(22635) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(22635))))  severity failure;
	assert RAM(22636) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22636))))  severity failure;
	assert RAM(22637) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(22637))))  severity failure;
	assert RAM(22638) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(22638))))  severity failure;
	assert RAM(22639) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(22639))))  severity failure;
	assert RAM(22640) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(22640))))  severity failure;
	assert RAM(22641) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22641))))  severity failure;
	assert RAM(22642) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(22642))))  severity failure;
	assert RAM(22643) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22643))))  severity failure;
	assert RAM(22644) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(22644))))  severity failure;
	assert RAM(22645) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(22645))))  severity failure;
	assert RAM(22646) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(22646))))  severity failure;
	assert RAM(22647) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(22647))))  severity failure;
	assert RAM(22648) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(22648))))  severity failure;
	assert RAM(22649) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22649))))  severity failure;
	assert RAM(22650) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(22650))))  severity failure;
	assert RAM(22651) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(22651))))  severity failure;
	assert RAM(22652) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(22652))))  severity failure;
	assert RAM(22653) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(22653))))  severity failure;
	assert RAM(22654) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(22654))))  severity failure;
	assert RAM(22655) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(22655))))  severity failure;
	assert RAM(22656) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(22656))))  severity failure;
	assert RAM(22657) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22657))))  severity failure;
	assert RAM(22658) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(22658))))  severity failure;
	assert RAM(22659) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(22659))))  severity failure;
	assert RAM(22660) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(22660))))  severity failure;
	assert RAM(22661) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22661))))  severity failure;
	assert RAM(22662) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(22662))))  severity failure;
	assert RAM(22663) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22663))))  severity failure;
	assert RAM(22664) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(22664))))  severity failure;
	assert RAM(22665) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22665))))  severity failure;
	assert RAM(22666) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(22666))))  severity failure;
	assert RAM(22667) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(22667))))  severity failure;
	assert RAM(22668) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(22668))))  severity failure;
	assert RAM(22669) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(22669))))  severity failure;
	assert RAM(22670) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22670))))  severity failure;
	assert RAM(22671) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(22671))))  severity failure;
	assert RAM(22672) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(22672))))  severity failure;
	assert RAM(22673) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(22673))))  severity failure;
	assert RAM(22674) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(22674))))  severity failure;
	assert RAM(22675) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(22675))))  severity failure;
	assert RAM(22676) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22676))))  severity failure;
	assert RAM(22677) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(22677))))  severity failure;
	assert RAM(22678) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(22678))))  severity failure;
	assert RAM(22679) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22679))))  severity failure;
	assert RAM(22680) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(22680))))  severity failure;
	assert RAM(22681) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(22681))))  severity failure;
	assert RAM(22682) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(22682))))  severity failure;
	assert RAM(22683) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(22683))))  severity failure;
	assert RAM(22684) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(22684))))  severity failure;
	assert RAM(22685) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(22685))))  severity failure;
	assert RAM(22686) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(22686))))  severity failure;
	assert RAM(22687) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22687))))  severity failure;
	assert RAM(22688) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(22688))))  severity failure;
	assert RAM(22689) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(22689))))  severity failure;
	assert RAM(22690) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(22690))))  severity failure;
	assert RAM(22691) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22691))))  severity failure;
	assert RAM(22692) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(22692))))  severity failure;
	assert RAM(22693) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(22693))))  severity failure;
	assert RAM(22694) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(22694))))  severity failure;
	assert RAM(22695) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(22695))))  severity failure;
	assert RAM(22696) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(22696))))  severity failure;
	assert RAM(22697) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(22697))))  severity failure;
	assert RAM(22698) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(22698))))  severity failure;
	assert RAM(22699) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(22699))))  severity failure;
	assert RAM(22700) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(22700))))  severity failure;
	assert RAM(22701) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(22701))))  severity failure;
	assert RAM(22702) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(22702))))  severity failure;
	assert RAM(22703) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(22703))))  severity failure;
	assert RAM(22704) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(22704))))  severity failure;
	assert RAM(22705) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(22705))))  severity failure;
	assert RAM(22706) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(22706))))  severity failure;
	assert RAM(22707) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(22707))))  severity failure;
	assert RAM(22708) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(22708))))  severity failure;
	assert RAM(22709) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(22709))))  severity failure;
	assert RAM(22710) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(22710))))  severity failure;
	assert RAM(22711) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(22711))))  severity failure;
	assert RAM(22712) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(22712))))  severity failure;
	assert RAM(22713) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22713))))  severity failure;
	assert RAM(22714) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(22714))))  severity failure;
	assert RAM(22715) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(22715))))  severity failure;
	assert RAM(22716) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(22716))))  severity failure;
	assert RAM(22717) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(22717))))  severity failure;
	assert RAM(22718) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22718))))  severity failure;
	assert RAM(22719) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(22719))))  severity failure;
	assert RAM(22720) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22720))))  severity failure;
	assert RAM(22721) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(22721))))  severity failure;
	assert RAM(22722) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(22722))))  severity failure;
	assert RAM(22723) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(22723))))  severity failure;
	assert RAM(22724) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(22724))))  severity failure;
	assert RAM(22725) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(22725))))  severity failure;
	assert RAM(22726) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22726))))  severity failure;
	assert RAM(22727) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(22727))))  severity failure;
	assert RAM(22728) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(22728))))  severity failure;
	assert RAM(22729) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(22729))))  severity failure;
	assert RAM(22730) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(22730))))  severity failure;
	assert RAM(22731) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22731))))  severity failure;
	assert RAM(22732) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(22732))))  severity failure;
	assert RAM(22733) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(22733))))  severity failure;
	assert RAM(22734) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(22734))))  severity failure;
	assert RAM(22735) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(22735))))  severity failure;
	assert RAM(22736) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(22736))))  severity failure;
	assert RAM(22737) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(22737))))  severity failure;
	assert RAM(22738) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(22738))))  severity failure;
	assert RAM(22739) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(22739))))  severity failure;
	assert RAM(22740) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(22740))))  severity failure;
	assert RAM(22741) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(22741))))  severity failure;
	assert RAM(22742) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(22742))))  severity failure;
	assert RAM(22743) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22743))))  severity failure;
	assert RAM(22744) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22744))))  severity failure;
	assert RAM(22745) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22745))))  severity failure;
	assert RAM(22746) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(22746))))  severity failure;
	assert RAM(22747) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(22747))))  severity failure;
	assert RAM(22748) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(22748))))  severity failure;
	assert RAM(22749) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(22749))))  severity failure;
	assert RAM(22750) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(22750))))  severity failure;
	assert RAM(22751) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(22751))))  severity failure;
	assert RAM(22752) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(22752))))  severity failure;
	assert RAM(22753) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(22753))))  severity failure;
	assert RAM(22754) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(22754))))  severity failure;
	assert RAM(22755) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(22755))))  severity failure;
	assert RAM(22756) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(22756))))  severity failure;
	assert RAM(22757) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(22757))))  severity failure;
	assert RAM(22758) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(22758))))  severity failure;
	assert RAM(22759) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(22759))))  severity failure;
	assert RAM(22760) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22760))))  severity failure;
	assert RAM(22761) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(22761))))  severity failure;
	assert RAM(22762) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(22762))))  severity failure;
	assert RAM(22763) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(22763))))  severity failure;
	assert RAM(22764) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(22764))))  severity failure;
	assert RAM(22765) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(22765))))  severity failure;
	assert RAM(22766) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(22766))))  severity failure;
	assert RAM(22767) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(22767))))  severity failure;
	assert RAM(22768) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(22768))))  severity failure;
	assert RAM(22769) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(22769))))  severity failure;
	assert RAM(22770) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(22770))))  severity failure;
	assert RAM(22771) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(22771))))  severity failure;
	assert RAM(22772) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(22772))))  severity failure;
	assert RAM(22773) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22773))))  severity failure;
	assert RAM(22774) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22774))))  severity failure;
	assert RAM(22775) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22775))))  severity failure;
	assert RAM(22776) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22776))))  severity failure;
	assert RAM(22777) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22777))))  severity failure;
	assert RAM(22778) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(22778))))  severity failure;
	assert RAM(22779) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22779))))  severity failure;
	assert RAM(22780) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(22780))))  severity failure;
	assert RAM(22781) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(22781))))  severity failure;
	assert RAM(22782) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(22782))))  severity failure;
	assert RAM(22783) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(22783))))  severity failure;
	assert RAM(22784) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(22784))))  severity failure;
	assert RAM(22785) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(22785))))  severity failure;
	assert RAM(22786) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(22786))))  severity failure;
	assert RAM(22787) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(22787))))  severity failure;
	assert RAM(22788) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22788))))  severity failure;
	assert RAM(22789) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(22789))))  severity failure;
	assert RAM(22790) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(22790))))  severity failure;
	assert RAM(22791) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(22791))))  severity failure;
	assert RAM(22792) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(22792))))  severity failure;
	assert RAM(22793) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(22793))))  severity failure;
	assert RAM(22794) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(22794))))  severity failure;
	assert RAM(22795) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(22795))))  severity failure;
	assert RAM(22796) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(22796))))  severity failure;
	assert RAM(22797) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(22797))))  severity failure;
	assert RAM(22798) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(22798))))  severity failure;
	assert RAM(22799) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(22799))))  severity failure;
	assert RAM(22800) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22800))))  severity failure;
	assert RAM(22801) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(22801))))  severity failure;
	assert RAM(22802) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22802))))  severity failure;
	assert RAM(22803) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(22803))))  severity failure;
	assert RAM(22804) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22804))))  severity failure;
	assert RAM(22805) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(22805))))  severity failure;
	assert RAM(22806) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(22806))))  severity failure;
	assert RAM(22807) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(22807))))  severity failure;
	assert RAM(22808) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22808))))  severity failure;
	assert RAM(22809) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(22809))))  severity failure;
	assert RAM(22810) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(22810))))  severity failure;
	assert RAM(22811) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22811))))  severity failure;
	assert RAM(22812) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22812))))  severity failure;
	assert RAM(22813) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(22813))))  severity failure;
	assert RAM(22814) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(22814))))  severity failure;
	assert RAM(22815) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(22815))))  severity failure;
	assert RAM(22816) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(22816))))  severity failure;
	assert RAM(22817) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(22817))))  severity failure;
	assert RAM(22818) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(22818))))  severity failure;
	assert RAM(22819) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(22819))))  severity failure;
	assert RAM(22820) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(22820))))  severity failure;
	assert RAM(22821) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(22821))))  severity failure;
	assert RAM(22822) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(22822))))  severity failure;
	assert RAM(22823) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(22823))))  severity failure;
	assert RAM(22824) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(22824))))  severity failure;
	assert RAM(22825) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(22825))))  severity failure;
	assert RAM(22826) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(22826))))  severity failure;
	assert RAM(22827) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22827))))  severity failure;
	assert RAM(22828) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(22828))))  severity failure;
	assert RAM(22829) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22829))))  severity failure;
	assert RAM(22830) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(22830))))  severity failure;
	assert RAM(22831) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(22831))))  severity failure;
	assert RAM(22832) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(22832))))  severity failure;
	assert RAM(22833) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(22833))))  severity failure;
	assert RAM(22834) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(22834))))  severity failure;
	assert RAM(22835) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(22835))))  severity failure;
	assert RAM(22836) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22836))))  severity failure;
	assert RAM(22837) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(22837))))  severity failure;
	assert RAM(22838) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22838))))  severity failure;
	assert RAM(22839) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22839))))  severity failure;
	assert RAM(22840) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(22840))))  severity failure;
	assert RAM(22841) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22841))))  severity failure;
	assert RAM(22842) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(22842))))  severity failure;
	assert RAM(22843) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(22843))))  severity failure;
	assert RAM(22844) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(22844))))  severity failure;
	assert RAM(22845) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(22845))))  severity failure;
	assert RAM(22846) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22846))))  severity failure;
	assert RAM(22847) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22847))))  severity failure;
	assert RAM(22848) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(22848))))  severity failure;
	assert RAM(22849) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(22849))))  severity failure;
	assert RAM(22850) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(22850))))  severity failure;
	assert RAM(22851) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(22851))))  severity failure;
	assert RAM(22852) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(22852))))  severity failure;
	assert RAM(22853) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(22853))))  severity failure;
	assert RAM(22854) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(22854))))  severity failure;
	assert RAM(22855) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(22855))))  severity failure;
	assert RAM(22856) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22856))))  severity failure;
	assert RAM(22857) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22857))))  severity failure;
	assert RAM(22858) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22858))))  severity failure;
	assert RAM(22859) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(22859))))  severity failure;
	assert RAM(22860) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(22860))))  severity failure;
	assert RAM(22861) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(22861))))  severity failure;
	assert RAM(22862) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22862))))  severity failure;
	assert RAM(22863) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(22863))))  severity failure;
	assert RAM(22864) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(22864))))  severity failure;
	assert RAM(22865) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(22865))))  severity failure;
	assert RAM(22866) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22866))))  severity failure;
	assert RAM(22867) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(22867))))  severity failure;
	assert RAM(22868) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(22868))))  severity failure;
	assert RAM(22869) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(22869))))  severity failure;
	assert RAM(22870) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(22870))))  severity failure;
	assert RAM(22871) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22871))))  severity failure;
	assert RAM(22872) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(22872))))  severity failure;
	assert RAM(22873) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(22873))))  severity failure;
	assert RAM(22874) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22874))))  severity failure;
	assert RAM(22875) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22875))))  severity failure;
	assert RAM(22876) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(22876))))  severity failure;
	assert RAM(22877) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(22877))))  severity failure;
	assert RAM(22878) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(22878))))  severity failure;
	assert RAM(22879) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22879))))  severity failure;
	assert RAM(22880) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(22880))))  severity failure;
	assert RAM(22881) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(22881))))  severity failure;
	assert RAM(22882) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(22882))))  severity failure;
	assert RAM(22883) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(22883))))  severity failure;
	assert RAM(22884) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(22884))))  severity failure;
	assert RAM(22885) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(22885))))  severity failure;
	assert RAM(22886) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(22886))))  severity failure;
	assert RAM(22887) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22887))))  severity failure;
	assert RAM(22888) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(22888))))  severity failure;
	assert RAM(22889) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(22889))))  severity failure;
	assert RAM(22890) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(22890))))  severity failure;
	assert RAM(22891) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(22891))))  severity failure;
	assert RAM(22892) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(22892))))  severity failure;
	assert RAM(22893) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(22893))))  severity failure;
	assert RAM(22894) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(22894))))  severity failure;
	assert RAM(22895) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22895))))  severity failure;
	assert RAM(22896) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(22896))))  severity failure;
	assert RAM(22897) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(22897))))  severity failure;
	assert RAM(22898) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(22898))))  severity failure;
	assert RAM(22899) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22899))))  severity failure;
	assert RAM(22900) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(22900))))  severity failure;
	assert RAM(22901) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(22901))))  severity failure;
	assert RAM(22902) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(22902))))  severity failure;
	assert RAM(22903) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(22903))))  severity failure;
	assert RAM(22904) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(22904))))  severity failure;
	assert RAM(22905) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(22905))))  severity failure;
	assert RAM(22906) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(22906))))  severity failure;
	assert RAM(22907) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22907))))  severity failure;
	assert RAM(22908) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(22908))))  severity failure;
	assert RAM(22909) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(22909))))  severity failure;
	assert RAM(22910) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(22910))))  severity failure;
	assert RAM(22911) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(22911))))  severity failure;
	assert RAM(22912) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22912))))  severity failure;
	assert RAM(22913) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(22913))))  severity failure;
	assert RAM(22914) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(22914))))  severity failure;
	assert RAM(22915) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(22915))))  severity failure;
	assert RAM(22916) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22916))))  severity failure;
	assert RAM(22917) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(22917))))  severity failure;
	assert RAM(22918) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(22918))))  severity failure;
	assert RAM(22919) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(22919))))  severity failure;
	assert RAM(22920) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(22920))))  severity failure;
	assert RAM(22921) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(22921))))  severity failure;
	assert RAM(22922) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(22922))))  severity failure;
	assert RAM(22923) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(22923))))  severity failure;
	assert RAM(22924) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(22924))))  severity failure;
	assert RAM(22925) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(22925))))  severity failure;
	assert RAM(22926) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22926))))  severity failure;
	assert RAM(22927) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(22927))))  severity failure;
	assert RAM(22928) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(22928))))  severity failure;
	assert RAM(22929) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(22929))))  severity failure;
	assert RAM(22930) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(22930))))  severity failure;
	assert RAM(22931) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(22931))))  severity failure;
	assert RAM(22932) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(22932))))  severity failure;
	assert RAM(22933) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(22933))))  severity failure;
	assert RAM(22934) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(22934))))  severity failure;
	assert RAM(22935) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(22935))))  severity failure;
	assert RAM(22936) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(22936))))  severity failure;
	assert RAM(22937) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(22937))))  severity failure;
	assert RAM(22938) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(22938))))  severity failure;
	assert RAM(22939) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(22939))))  severity failure;
	assert RAM(22940) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(22940))))  severity failure;
	assert RAM(22941) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(22941))))  severity failure;
	assert RAM(22942) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(22942))))  severity failure;
	assert RAM(22943) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(22943))))  severity failure;
	assert RAM(22944) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(22944))))  severity failure;
	assert RAM(22945) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(22945))))  severity failure;
	assert RAM(22946) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(22946))))  severity failure;
	assert RAM(22947) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(22947))))  severity failure;
	assert RAM(22948) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(22948))))  severity failure;
	assert RAM(22949) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(22949))))  severity failure;
	assert RAM(22950) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(22950))))  severity failure;
	assert RAM(22951) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(22951))))  severity failure;
	assert RAM(22952) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(22952))))  severity failure;
	assert RAM(22953) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(22953))))  severity failure;
	assert RAM(22954) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(22954))))  severity failure;
	assert RAM(22955) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(22955))))  severity failure;
	assert RAM(22956) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(22956))))  severity failure;
	assert RAM(22957) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(22957))))  severity failure;
	assert RAM(22958) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(22958))))  severity failure;
	assert RAM(22959) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(22959))))  severity failure;
	assert RAM(22960) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(22960))))  severity failure;
	assert RAM(22961) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(22961))))  severity failure;
	assert RAM(22962) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(22962))))  severity failure;
	assert RAM(22963) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(22963))))  severity failure;
	assert RAM(22964) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(22964))))  severity failure;
	assert RAM(22965) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(22965))))  severity failure;
	assert RAM(22966) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(22966))))  severity failure;
	assert RAM(22967) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(22967))))  severity failure;
	assert RAM(22968) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(22968))))  severity failure;
	assert RAM(22969) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(22969))))  severity failure;
	assert RAM(22970) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(22970))))  severity failure;
	assert RAM(22971) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(22971))))  severity failure;
	assert RAM(22972) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(22972))))  severity failure;
	assert RAM(22973) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(22973))))  severity failure;
	assert RAM(22974) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(22974))))  severity failure;
	assert RAM(22975) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(22975))))  severity failure;
	assert RAM(22976) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(22976))))  severity failure;
	assert RAM(22977) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(22977))))  severity failure;
	assert RAM(22978) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(22978))))  severity failure;
	assert RAM(22979) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(22979))))  severity failure;
	assert RAM(22980) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(22980))))  severity failure;
	assert RAM(22981) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(22981))))  severity failure;
	assert RAM(22982) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(22982))))  severity failure;
	assert RAM(22983) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(22983))))  severity failure;
	assert RAM(22984) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(22984))))  severity failure;
	assert RAM(22985) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(22985))))  severity failure;
	assert RAM(22986) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(22986))))  severity failure;
	assert RAM(22987) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(22987))))  severity failure;
	assert RAM(22988) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22988))))  severity failure;
	assert RAM(22989) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(22989))))  severity failure;
	assert RAM(22990) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(22990))))  severity failure;
	assert RAM(22991) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(22991))))  severity failure;
	assert RAM(22992) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(22992))))  severity failure;
	assert RAM(22993) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(22993))))  severity failure;
	assert RAM(22994) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(22994))))  severity failure;
	assert RAM(22995) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(22995))))  severity failure;
	assert RAM(22996) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(22996))))  severity failure;
	assert RAM(22997) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(22997))))  severity failure;
	assert RAM(22998) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(22998))))  severity failure;
	assert RAM(22999) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(22999))))  severity failure;
	assert RAM(23000) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(23000))))  severity failure;
	assert RAM(23001) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(23001))))  severity failure;
	assert RAM(23002) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(23002))))  severity failure;
	assert RAM(23003) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(23003))))  severity failure;
	assert RAM(23004) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(23004))))  severity failure;
	assert RAM(23005) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(23005))))  severity failure;
	assert RAM(23006) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(23006))))  severity failure;
	assert RAM(23007) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(23007))))  severity failure;
	assert RAM(23008) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(23008))))  severity failure;
	assert RAM(23009) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(23009))))  severity failure;
	assert RAM(23010) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(23010))))  severity failure;
	assert RAM(23011) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(23011))))  severity failure;
	assert RAM(23012) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(23012))))  severity failure;
	assert RAM(23013) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(23013))))  severity failure;
	assert RAM(23014) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(23014))))  severity failure;
	assert RAM(23015) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(23015))))  severity failure;
	assert RAM(23016) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(23016))))  severity failure;
	assert RAM(23017) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(23017))))  severity failure;
	assert RAM(23018) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(23018))))  severity failure;
	assert RAM(23019) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(23019))))  severity failure;
	assert RAM(23020) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(23020))))  severity failure;
	assert RAM(23021) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(23021))))  severity failure;
	assert RAM(23022) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(23022))))  severity failure;
	assert RAM(23023) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(23023))))  severity failure;
	assert RAM(23024) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(23024))))  severity failure;
	assert RAM(23025) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(23025))))  severity failure;
	assert RAM(23026) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(23026))))  severity failure;
	assert RAM(23027) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(23027))))  severity failure;
	assert RAM(23028) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(23028))))  severity failure;
	assert RAM(23029) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(23029))))  severity failure;
	assert RAM(23030) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(23030))))  severity failure;
	assert RAM(23031) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(23031))))  severity failure;
	assert RAM(23032) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(23032))))  severity failure;
	assert RAM(23033) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(23033))))  severity failure;
	assert RAM(23034) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(23034))))  severity failure;
	assert RAM(23035) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(23035))))  severity failure;
	assert RAM(23036) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(23036))))  severity failure;
	assert RAM(23037) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(23037))))  severity failure;
	assert RAM(23038) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(23038))))  severity failure;
	assert RAM(23039) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(23039))))  severity failure;
	assert RAM(23040) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(23040))))  severity failure;
	assert RAM(23041) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(23041))))  severity failure;
	assert RAM(23042) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(23042))))  severity failure;
	assert RAM(23043) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(23043))))  severity failure;
	assert RAM(23044) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(23044))))  severity failure;
	assert RAM(23045) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(23045))))  severity failure;
	assert RAM(23046) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(23046))))  severity failure;
	assert RAM(23047) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(23047))))  severity failure;
	assert RAM(23048) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(23048))))  severity failure;
	assert RAM(23049) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(23049))))  severity failure;
	assert RAM(23050) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(23050))))  severity failure;
	assert RAM(23051) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(23051))))  severity failure;
	assert RAM(23052) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(23052))))  severity failure;
	assert RAM(23053) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(23053))))  severity failure;
	assert RAM(23054) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(23054))))  severity failure;
	assert RAM(23055) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(23055))))  severity failure;
	assert RAM(23056) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(23056))))  severity failure;
	assert RAM(23057) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(23057))))  severity failure;
	assert RAM(23058) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(23058))))  severity failure;
	assert RAM(23059) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(23059))))  severity failure;
	assert RAM(23060) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(23060))))  severity failure;
	assert RAM(23061) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(23061))))  severity failure;
	assert RAM(23062) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(23062))))  severity failure;
	assert RAM(23063) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(23063))))  severity failure;
	assert RAM(23064) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(23064))))  severity failure;
	assert RAM(23065) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(23065))))  severity failure;
	assert RAM(23066) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(23066))))  severity failure;
	assert RAM(23067) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(23067))))  severity failure;
	assert RAM(23068) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(23068))))  severity failure;
	assert RAM(23069) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(23069))))  severity failure;
	assert RAM(23070) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(23070))))  severity failure;
	assert RAM(23071) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(23071))))  severity failure;
	assert RAM(23072) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(23072))))  severity failure;
	assert RAM(23073) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(23073))))  severity failure;
	assert RAM(23074) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(23074))))  severity failure;
	assert RAM(23075) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(23075))))  severity failure;
	assert RAM(23076) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(23076))))  severity failure;
	assert RAM(23077) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23077))))  severity failure;
	assert RAM(23078) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(23078))))  severity failure;
	assert RAM(23079) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(23079))))  severity failure;
	assert RAM(23080) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(23080))))  severity failure;
	assert RAM(23081) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(23081))))  severity failure;
	assert RAM(23082) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(23082))))  severity failure;
	assert RAM(23083) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(23083))))  severity failure;
	assert RAM(23084) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(23084))))  severity failure;
	assert RAM(23085) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(23085))))  severity failure;
	assert RAM(23086) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(23086))))  severity failure;
	assert RAM(23087) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(23087))))  severity failure;
	assert RAM(23088) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(23088))))  severity failure;
	assert RAM(23089) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(23089))))  severity failure;
	assert RAM(23090) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(23090))))  severity failure;
	assert RAM(23091) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(23091))))  severity failure;
	assert RAM(23092) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(23092))))  severity failure;
	assert RAM(23093) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(23093))))  severity failure;
	assert RAM(23094) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(23094))))  severity failure;
	assert RAM(23095) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(23095))))  severity failure;
	assert RAM(23096) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(23096))))  severity failure;
	assert RAM(23097) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(23097))))  severity failure;
	assert RAM(23098) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(23098))))  severity failure;
	assert RAM(23099) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(23099))))  severity failure;
	assert RAM(23100) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(23100))))  severity failure;
	assert RAM(23101) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(23101))))  severity failure;
	assert RAM(23102) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(23102))))  severity failure;
	assert RAM(23103) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(23103))))  severity failure;
	assert RAM(23104) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(23104))))  severity failure;
	assert RAM(23105) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(23105))))  severity failure;
	assert RAM(23106) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(23106))))  severity failure;
	assert RAM(23107) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(23107))))  severity failure;
	assert RAM(23108) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(23108))))  severity failure;
	assert RAM(23109) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(23109))))  severity failure;
	assert RAM(23110) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(23110))))  severity failure;
	assert RAM(23111) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(23111))))  severity failure;
	assert RAM(23112) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(23112))))  severity failure;
	assert RAM(23113) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(23113))))  severity failure;
	assert RAM(23114) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(23114))))  severity failure;
	assert RAM(23115) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(23115))))  severity failure;
	assert RAM(23116) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(23116))))  severity failure;
	assert RAM(23117) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(23117))))  severity failure;
	assert RAM(23118) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(23118))))  severity failure;
	assert RAM(23119) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(23119))))  severity failure;
	assert RAM(23120) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(23120))))  severity failure;
	assert RAM(23121) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(23121))))  severity failure;
	assert RAM(23122) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(23122))))  severity failure;
	assert RAM(23123) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(23123))))  severity failure;
	assert RAM(23124) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(23124))))  severity failure;
	assert RAM(23125) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(23125))))  severity failure;
	assert RAM(23126) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(23126))))  severity failure;
	assert RAM(23127) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(23127))))  severity failure;
	assert RAM(23128) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(23128))))  severity failure;
	assert RAM(23129) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(23129))))  severity failure;
	assert RAM(23130) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(23130))))  severity failure;
	assert RAM(23131) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(23131))))  severity failure;
	assert RAM(23132) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(23132))))  severity failure;
	assert RAM(23133) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(23133))))  severity failure;
	assert RAM(23134) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(23134))))  severity failure;
	assert RAM(23135) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(23135))))  severity failure;
	assert RAM(23136) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(23136))))  severity failure;
	assert RAM(23137) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(23137))))  severity failure;
	assert RAM(23138) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(23138))))  severity failure;
	assert RAM(23139) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(23139))))  severity failure;
	assert RAM(23140) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(23140))))  severity failure;
	assert RAM(23141) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(23141))))  severity failure;
	assert RAM(23142) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(23142))))  severity failure;
	assert RAM(23143) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(23143))))  severity failure;
	assert RAM(23144) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(23144))))  severity failure;
	assert RAM(23145) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(23145))))  severity failure;
	assert RAM(23146) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(23146))))  severity failure;
	assert RAM(23147) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(23147))))  severity failure;
	assert RAM(23148) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(23148))))  severity failure;
	assert RAM(23149) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(23149))))  severity failure;
	assert RAM(23150) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(23150))))  severity failure;
	assert RAM(23151) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(23151))))  severity failure;
	assert RAM(23152) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(23152))))  severity failure;
	assert RAM(23153) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(23153))))  severity failure;
	assert RAM(23154) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(23154))))  severity failure;
	assert RAM(23155) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(23155))))  severity failure;
	assert RAM(23156) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(23156))))  severity failure;
	assert RAM(23157) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(23157))))  severity failure;
	assert RAM(23158) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(23158))))  severity failure;
	assert RAM(23159) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(23159))))  severity failure;
	assert RAM(23160) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(23160))))  severity failure;
	assert RAM(23161) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(23161))))  severity failure;
	assert RAM(23162) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(23162))))  severity failure;
	assert RAM(23163) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(23163))))  severity failure;
	assert RAM(23164) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(23164))))  severity failure;
	assert RAM(23165) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(23165))))  severity failure;
	assert RAM(23166) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(23166))))  severity failure;
	assert RAM(23167) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(23167))))  severity failure;
	assert RAM(23168) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(23168))))  severity failure;
	assert RAM(23169) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(23169))))  severity failure;
	assert RAM(23170) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(23170))))  severity failure;
	assert RAM(23171) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(23171))))  severity failure;
	assert RAM(23172) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(23172))))  severity failure;
	assert RAM(23173) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(23173))))  severity failure;
	assert RAM(23174) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(23174))))  severity failure;
	assert RAM(23175) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(23175))))  severity failure;
	assert RAM(23176) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(23176))))  severity failure;
	assert RAM(23177) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(23177))))  severity failure;
	assert RAM(23178) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(23178))))  severity failure;
	assert RAM(23179) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(23179))))  severity failure;
	assert RAM(23180) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(23180))))  severity failure;
	assert RAM(23181) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(23181))))  severity failure;
	assert RAM(23182) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(23182))))  severity failure;
	assert RAM(23183) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(23183))))  severity failure;
	assert RAM(23184) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(23184))))  severity failure;
	assert RAM(23185) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(23185))))  severity failure;
	assert RAM(23186) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(23186))))  severity failure;
	assert RAM(23187) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(23187))))  severity failure;
	assert RAM(23188) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(23188))))  severity failure;
	assert RAM(23189) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(23189))))  severity failure;
	assert RAM(23190) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(23190))))  severity failure;
	assert RAM(23191) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(23191))))  severity failure;
	assert RAM(23192) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(23192))))  severity failure;
	assert RAM(23193) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(23193))))  severity failure;
	assert RAM(23194) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(23194))))  severity failure;
	assert RAM(23195) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(23195))))  severity failure;
	assert RAM(23196) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(23196))))  severity failure;
	assert RAM(23197) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(23197))))  severity failure;
	assert RAM(23198) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(23198))))  severity failure;
	assert RAM(23199) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(23199))))  severity failure;
	assert RAM(23200) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(23200))))  severity failure;
	assert RAM(23201) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(23201))))  severity failure;
	assert RAM(23202) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(23202))))  severity failure;
	assert RAM(23203) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(23203))))  severity failure;
	assert RAM(23204) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(23204))))  severity failure;
	assert RAM(23205) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(23205))))  severity failure;
	assert RAM(23206) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(23206))))  severity failure;
	assert RAM(23207) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(23207))))  severity failure;
	assert RAM(23208) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(23208))))  severity failure;
	assert RAM(23209) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(23209))))  severity failure;
	assert RAM(23210) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(23210))))  severity failure;
	assert RAM(23211) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(23211))))  severity failure;
	assert RAM(23212) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(23212))))  severity failure;
	assert RAM(23213) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(23213))))  severity failure;
	assert RAM(23214) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(23214))))  severity failure;
	assert RAM(23215) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(23215))))  severity failure;
	assert RAM(23216) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(23216))))  severity failure;
	assert RAM(23217) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(23217))))  severity failure;
	assert RAM(23218) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(23218))))  severity failure;
	assert RAM(23219) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(23219))))  severity failure;
	assert RAM(23220) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(23220))))  severity failure;
	assert RAM(23221) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(23221))))  severity failure;
	assert RAM(23222) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(23222))))  severity failure;
	assert RAM(23223) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(23223))))  severity failure;
	assert RAM(23224) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(23224))))  severity failure;
	assert RAM(23225) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(23225))))  severity failure;
	assert RAM(23226) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(23226))))  severity failure;
	assert RAM(23227) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(23227))))  severity failure;
	assert RAM(23228) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(23228))))  severity failure;
	assert RAM(23229) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(23229))))  severity failure;
	assert RAM(23230) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(23230))))  severity failure;
	assert RAM(23231) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(23231))))  severity failure;
	assert RAM(23232) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(23232))))  severity failure;
	assert RAM(23233) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(23233))))  severity failure;
	assert RAM(23234) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(23234))))  severity failure;
	assert RAM(23235) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(23235))))  severity failure;
	assert RAM(23236) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(23236))))  severity failure;
	assert RAM(23237) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(23237))))  severity failure;
	assert RAM(23238) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(23238))))  severity failure;
	assert RAM(23239) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(23239))))  severity failure;
	assert RAM(23240) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(23240))))  severity failure;
	assert RAM(23241) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(23241))))  severity failure;
	assert RAM(23242) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(23242))))  severity failure;
	assert RAM(23243) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(23243))))  severity failure;
	assert RAM(23244) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(23244))))  severity failure;
	assert RAM(23245) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(23245))))  severity failure;
	assert RAM(23246) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(23246))))  severity failure;
	assert RAM(23247) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(23247))))  severity failure;
	assert RAM(23248) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(23248))))  severity failure;
	assert RAM(23249) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(23249))))  severity failure;
	assert RAM(23250) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(23250))))  severity failure;
	assert RAM(23251) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(23251))))  severity failure;
	assert RAM(23252) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(23252))))  severity failure;
	assert RAM(23253) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(23253))))  severity failure;
	assert RAM(23254) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(23254))))  severity failure;
	assert RAM(23255) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(23255))))  severity failure;
	assert RAM(23256) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(23256))))  severity failure;
	assert RAM(23257) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(23257))))  severity failure;
	assert RAM(23258) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(23258))))  severity failure;
	assert RAM(23259) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(23259))))  severity failure;
	assert RAM(23260) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(23260))))  severity failure;
	assert RAM(23261) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(23261))))  severity failure;
	assert RAM(23262) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(23262))))  severity failure;
	assert RAM(23263) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(23263))))  severity failure;
	assert RAM(23264) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(23264))))  severity failure;
	assert RAM(23265) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(23265))))  severity failure;
	assert RAM(23266) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(23266))))  severity failure;
	assert RAM(23267) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(23267))))  severity failure;
	assert RAM(23268) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(23268))))  severity failure;
	assert RAM(23269) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(23269))))  severity failure;
	assert RAM(23270) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(23270))))  severity failure;
	assert RAM(23271) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(23271))))  severity failure;
	assert RAM(23272) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(23272))))  severity failure;
	assert RAM(23273) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(23273))))  severity failure;
	assert RAM(23274) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(23274))))  severity failure;
	assert RAM(23275) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(23275))))  severity failure;
	assert RAM(23276) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(23276))))  severity failure;
	assert RAM(23277) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(23277))))  severity failure;
	assert RAM(23278) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(23278))))  severity failure;
	assert RAM(23279) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(23279))))  severity failure;
	assert RAM(23280) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(23280))))  severity failure;
	assert RAM(23281) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(23281))))  severity failure;
    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;
end projecttb;
