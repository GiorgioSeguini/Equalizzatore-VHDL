library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
entity project_tb is
end project_tb;
architecture projecttb of project_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;
type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (
			0 => std_logic_vector(to_unsigned(27, 8)),
			1 => std_logic_vector(to_unsigned(90, 8)),
			2 => std_logic_vector(to_unsigned(224, 8)),
			3 => std_logic_vector(to_unsigned(113, 8)),
			4 => std_logic_vector(to_unsigned(53, 8)),
			5 => std_logic_vector(to_unsigned(100, 8)),
			6 => std_logic_vector(to_unsigned(63, 8)),
			7 => std_logic_vector(to_unsigned(138, 8)),
			8 => std_logic_vector(to_unsigned(207, 8)),
			9 => std_logic_vector(to_unsigned(199, 8)),
			10 => std_logic_vector(to_unsigned(222, 8)),
			11 => std_logic_vector(to_unsigned(149, 8)),
			12 => std_logic_vector(to_unsigned(39, 8)),
			13 => std_logic_vector(to_unsigned(221, 8)),
			14 => std_logic_vector(to_unsigned(231, 8)),
			15 => std_logic_vector(to_unsigned(103, 8)),
			16 => std_logic_vector(to_unsigned(217, 8)),
			17 => std_logic_vector(to_unsigned(252, 8)),
			18 => std_logic_vector(to_unsigned(53, 8)),
			19 => std_logic_vector(to_unsigned(211, 8)),
			20 => std_logic_vector(to_unsigned(243, 8)),
			21 => std_logic_vector(to_unsigned(213, 8)),
			22 => std_logic_vector(to_unsigned(150, 8)),
			23 => std_logic_vector(to_unsigned(157, 8)),
			24 => std_logic_vector(to_unsigned(128, 8)),
			25 => std_logic_vector(to_unsigned(31, 8)),
			26 => std_logic_vector(to_unsigned(171, 8)),
			27 => std_logic_vector(to_unsigned(209, 8)),
			28 => std_logic_vector(to_unsigned(24, 8)),
			29 => std_logic_vector(to_unsigned(148, 8)),
			30 => std_logic_vector(to_unsigned(4, 8)),
			31 => std_logic_vector(to_unsigned(106, 8)),
			32 => std_logic_vector(to_unsigned(138, 8)),
			33 => std_logic_vector(to_unsigned(171, 8)),
			34 => std_logic_vector(to_unsigned(103, 8)),
			35 => std_logic_vector(to_unsigned(26, 8)),
			36 => std_logic_vector(to_unsigned(90, 8)),
			37 => std_logic_vector(to_unsigned(2, 8)),
			38 => std_logic_vector(to_unsigned(21, 8)),
			39 => std_logic_vector(to_unsigned(23, 8)),
			40 => std_logic_vector(to_unsigned(169, 8)),
			41 => std_logic_vector(to_unsigned(196, 8)),
			42 => std_logic_vector(to_unsigned(151, 8)),
			43 => std_logic_vector(to_unsigned(193, 8)),
			44 => std_logic_vector(to_unsigned(255, 8)),
			45 => std_logic_vector(to_unsigned(229, 8)),
			46 => std_logic_vector(to_unsigned(138, 8)),
			47 => std_logic_vector(to_unsigned(47, 8)),
			48 => std_logic_vector(to_unsigned(58, 8)),
			49 => std_logic_vector(to_unsigned(223, 8)),
			50 => std_logic_vector(to_unsigned(54, 8)),
			51 => std_logic_vector(to_unsigned(82, 8)),
			52 => std_logic_vector(to_unsigned(222, 8)),
			53 => std_logic_vector(to_unsigned(101, 8)),
			54 => std_logic_vector(to_unsigned(226, 8)),
			55 => std_logic_vector(to_unsigned(146, 8)),
			56 => std_logic_vector(to_unsigned(67, 8)),
			57 => std_logic_vector(to_unsigned(106, 8)),
			58 => std_logic_vector(to_unsigned(11, 8)),
			59 => std_logic_vector(to_unsigned(10, 8)),
			60 => std_logic_vector(to_unsigned(65, 8)),
			61 => std_logic_vector(to_unsigned(189, 8)),
			62 => std_logic_vector(to_unsigned(118, 8)),
			63 => std_logic_vector(to_unsigned(14, 8)),
			64 => std_logic_vector(to_unsigned(151, 8)),
			65 => std_logic_vector(to_unsigned(139, 8)),
			66 => std_logic_vector(to_unsigned(3, 8)),
			67 => std_logic_vector(to_unsigned(134, 8)),
			68 => std_logic_vector(to_unsigned(221, 8)),
			69 => std_logic_vector(to_unsigned(229, 8)),
			70 => std_logic_vector(to_unsigned(235, 8)),
			71 => std_logic_vector(to_unsigned(188, 8)),
			72 => std_logic_vector(to_unsigned(27, 8)),
			73 => std_logic_vector(to_unsigned(171, 8)),
			74 => std_logic_vector(to_unsigned(248, 8)),
			75 => std_logic_vector(to_unsigned(139, 8)),
			76 => std_logic_vector(to_unsigned(111, 8)),
			77 => std_logic_vector(to_unsigned(82, 8)),
			78 => std_logic_vector(to_unsigned(254, 8)),
			79 => std_logic_vector(to_unsigned(31, 8)),
			80 => std_logic_vector(to_unsigned(127, 8)),
			81 => std_logic_vector(to_unsigned(193, 8)),
			82 => std_logic_vector(to_unsigned(182, 8)),
			83 => std_logic_vector(to_unsigned(136, 8)),
			84 => std_logic_vector(to_unsigned(74, 8)),
			85 => std_logic_vector(to_unsigned(217, 8)),
			86 => std_logic_vector(to_unsigned(184, 8)),
			87 => std_logic_vector(to_unsigned(186, 8)),
			88 => std_logic_vector(to_unsigned(41, 8)),
			89 => std_logic_vector(to_unsigned(185, 8)),
			90 => std_logic_vector(to_unsigned(232, 8)),
			91 => std_logic_vector(to_unsigned(98, 8)),
			92 => std_logic_vector(to_unsigned(229, 8)),
			93 => std_logic_vector(to_unsigned(236, 8)),
			94 => std_logic_vector(to_unsigned(250, 8)),
			95 => std_logic_vector(to_unsigned(118, 8)),
			96 => std_logic_vector(to_unsigned(252, 8)),
			97 => std_logic_vector(to_unsigned(66, 8)),
			98 => std_logic_vector(to_unsigned(116, 8)),
			99 => std_logic_vector(to_unsigned(37, 8)),
			100 => std_logic_vector(to_unsigned(248, 8)),
			101 => std_logic_vector(to_unsigned(22, 8)),
			102 => std_logic_vector(to_unsigned(38, 8)),
			103 => std_logic_vector(to_unsigned(75, 8)),
			104 => std_logic_vector(to_unsigned(207, 8)),
			105 => std_logic_vector(to_unsigned(14, 8)),
			106 => std_logic_vector(to_unsigned(123, 8)),
			107 => std_logic_vector(to_unsigned(32, 8)),
			108 => std_logic_vector(to_unsigned(200, 8)),
			109 => std_logic_vector(to_unsigned(171, 8)),
			110 => std_logic_vector(to_unsigned(150, 8)),
			111 => std_logic_vector(to_unsigned(76, 8)),
			112 => std_logic_vector(to_unsigned(112, 8)),
			113 => std_logic_vector(to_unsigned(254, 8)),
			114 => std_logic_vector(to_unsigned(73, 8)),
			115 => std_logic_vector(to_unsigned(70, 8)),
			116 => std_logic_vector(to_unsigned(26, 8)),
			117 => std_logic_vector(to_unsigned(56, 8)),
			118 => std_logic_vector(to_unsigned(151, 8)),
			119 => std_logic_vector(to_unsigned(196, 8)),
			120 => std_logic_vector(to_unsigned(248, 8)),
			121 => std_logic_vector(to_unsigned(196, 8)),
			122 => std_logic_vector(to_unsigned(182, 8)),
			123 => std_logic_vector(to_unsigned(163, 8)),
			124 => std_logic_vector(to_unsigned(32, 8)),
			125 => std_logic_vector(to_unsigned(35, 8)),
			126 => std_logic_vector(to_unsigned(8, 8)),
			127 => std_logic_vector(to_unsigned(119, 8)),
			128 => std_logic_vector(to_unsigned(193, 8)),
			129 => std_logic_vector(to_unsigned(81, 8)),
			130 => std_logic_vector(to_unsigned(22, 8)),
			131 => std_logic_vector(to_unsigned(157, 8)),
			132 => std_logic_vector(to_unsigned(217, 8)),
			133 => std_logic_vector(to_unsigned(128, 8)),
			134 => std_logic_vector(to_unsigned(76, 8)),
			135 => std_logic_vector(to_unsigned(143, 8)),
			136 => std_logic_vector(to_unsigned(188, 8)),
			137 => std_logic_vector(to_unsigned(73, 8)),
			138 => std_logic_vector(to_unsigned(239, 8)),
			139 => std_logic_vector(to_unsigned(83, 8)),
			140 => std_logic_vector(to_unsigned(129, 8)),
			141 => std_logic_vector(to_unsigned(145, 8)),
			142 => std_logic_vector(to_unsigned(217, 8)),
			143 => std_logic_vector(to_unsigned(11, 8)),
			144 => std_logic_vector(to_unsigned(183, 8)),
			145 => std_logic_vector(to_unsigned(254, 8)),
			146 => std_logic_vector(to_unsigned(30, 8)),
			147 => std_logic_vector(to_unsigned(18, 8)),
			148 => std_logic_vector(to_unsigned(223, 8)),
			149 => std_logic_vector(to_unsigned(1, 8)),
			150 => std_logic_vector(to_unsigned(107, 8)),
			151 => std_logic_vector(to_unsigned(126, 8)),
			152 => std_logic_vector(to_unsigned(44, 8)),
			153 => std_logic_vector(to_unsigned(73, 8)),
			154 => std_logic_vector(to_unsigned(211, 8)),
			155 => std_logic_vector(to_unsigned(151, 8)),
			156 => std_logic_vector(to_unsigned(145, 8)),
			157 => std_logic_vector(to_unsigned(156, 8)),
			158 => std_logic_vector(to_unsigned(252, 8)),
			159 => std_logic_vector(to_unsigned(27, 8)),
			160 => std_logic_vector(to_unsigned(7, 8)),
			161 => std_logic_vector(to_unsigned(146, 8)),
			162 => std_logic_vector(to_unsigned(206, 8)),
			163 => std_logic_vector(to_unsigned(71, 8)),
			164 => std_logic_vector(to_unsigned(173, 8)),
			165 => std_logic_vector(to_unsigned(72, 8)),
			166 => std_logic_vector(to_unsigned(65, 8)),
			167 => std_logic_vector(to_unsigned(69, 8)),
			168 => std_logic_vector(to_unsigned(205, 8)),
			169 => std_logic_vector(to_unsigned(119, 8)),
			170 => std_logic_vector(to_unsigned(43, 8)),
			171 => std_logic_vector(to_unsigned(189, 8)),
			172 => std_logic_vector(to_unsigned(92, 8)),
			173 => std_logic_vector(to_unsigned(243, 8)),
			174 => std_logic_vector(to_unsigned(20, 8)),
			175 => std_logic_vector(to_unsigned(111, 8)),
			176 => std_logic_vector(to_unsigned(64, 8)),
			177 => std_logic_vector(to_unsigned(179, 8)),
			178 => std_logic_vector(to_unsigned(88, 8)),
			179 => std_logic_vector(to_unsigned(151, 8)),
			180 => std_logic_vector(to_unsigned(209, 8)),
			181 => std_logic_vector(to_unsigned(87, 8)),
			182 => std_logic_vector(to_unsigned(220, 8)),
			183 => std_logic_vector(to_unsigned(34, 8)),
			184 => std_logic_vector(to_unsigned(196, 8)),
			185 => std_logic_vector(to_unsigned(199, 8)),
			186 => std_logic_vector(to_unsigned(205, 8)),
			187 => std_logic_vector(to_unsigned(83, 8)),
			188 => std_logic_vector(to_unsigned(88, 8)),
			189 => std_logic_vector(to_unsigned(123, 8)),
			190 => std_logic_vector(to_unsigned(69, 8)),
			191 => std_logic_vector(to_unsigned(219, 8)),
			192 => std_logic_vector(to_unsigned(57, 8)),
			193 => std_logic_vector(to_unsigned(165, 8)),
			194 => std_logic_vector(to_unsigned(34, 8)),
			195 => std_logic_vector(to_unsigned(242, 8)),
			196 => std_logic_vector(to_unsigned(180, 8)),
			197 => std_logic_vector(to_unsigned(238, 8)),
			198 => std_logic_vector(to_unsigned(105, 8)),
			199 => std_logic_vector(to_unsigned(176, 8)),
			200 => std_logic_vector(to_unsigned(217, 8)),
			201 => std_logic_vector(to_unsigned(84, 8)),
			202 => std_logic_vector(to_unsigned(9, 8)),
			203 => std_logic_vector(to_unsigned(247, 8)),
			204 => std_logic_vector(to_unsigned(95, 8)),
			205 => std_logic_vector(to_unsigned(35, 8)),
			206 => std_logic_vector(to_unsigned(193, 8)),
			207 => std_logic_vector(to_unsigned(125, 8)),
			208 => std_logic_vector(to_unsigned(131, 8)),
			209 => std_logic_vector(to_unsigned(142, 8)),
			210 => std_logic_vector(to_unsigned(205, 8)),
			211 => std_logic_vector(to_unsigned(201, 8)),
			212 => std_logic_vector(to_unsigned(135, 8)),
			213 => std_logic_vector(to_unsigned(84, 8)),
			214 => std_logic_vector(to_unsigned(187, 8)),
			215 => std_logic_vector(to_unsigned(138, 8)),
			216 => std_logic_vector(to_unsigned(116, 8)),
			217 => std_logic_vector(to_unsigned(94, 8)),
			218 => std_logic_vector(to_unsigned(121, 8)),
			219 => std_logic_vector(to_unsigned(149, 8)),
			220 => std_logic_vector(to_unsigned(73, 8)),
			221 => std_logic_vector(to_unsigned(121, 8)),
			222 => std_logic_vector(to_unsigned(160, 8)),
			223 => std_logic_vector(to_unsigned(120, 8)),
			224 => std_logic_vector(to_unsigned(137, 8)),
			225 => std_logic_vector(to_unsigned(136, 8)),
			226 => std_logic_vector(to_unsigned(249, 8)),
			227 => std_logic_vector(to_unsigned(201, 8)),
			228 => std_logic_vector(to_unsigned(111, 8)),
			229 => std_logic_vector(to_unsigned(210, 8)),
			230 => std_logic_vector(to_unsigned(140, 8)),
			231 => std_logic_vector(to_unsigned(95, 8)),
			232 => std_logic_vector(to_unsigned(170, 8)),
			233 => std_logic_vector(to_unsigned(65, 8)),
			234 => std_logic_vector(to_unsigned(230, 8)),
			235 => std_logic_vector(to_unsigned(129, 8)),
			236 => std_logic_vector(to_unsigned(152, 8)),
			237 => std_logic_vector(to_unsigned(240, 8)),
			238 => std_logic_vector(to_unsigned(149, 8)),
			239 => std_logic_vector(to_unsigned(192, 8)),
			240 => std_logic_vector(to_unsigned(85, 8)),
			241 => std_logic_vector(to_unsigned(211, 8)),
			242 => std_logic_vector(to_unsigned(128, 8)),
			243 => std_logic_vector(to_unsigned(32, 8)),
			244 => std_logic_vector(to_unsigned(38, 8)),
			245 => std_logic_vector(to_unsigned(78, 8)),
			246 => std_logic_vector(to_unsigned(235, 8)),
			247 => std_logic_vector(to_unsigned(108, 8)),
			248 => std_logic_vector(to_unsigned(125, 8)),
			249 => std_logic_vector(to_unsigned(100, 8)),
			250 => std_logic_vector(to_unsigned(87, 8)),
			251 => std_logic_vector(to_unsigned(10, 8)),
			252 => std_logic_vector(to_unsigned(238, 8)),
			253 => std_logic_vector(to_unsigned(197, 8)),
			254 => std_logic_vector(to_unsigned(185, 8)),
			255 => std_logic_vector(to_unsigned(244, 8)),
			256 => std_logic_vector(to_unsigned(228, 8)),
			257 => std_logic_vector(to_unsigned(81, 8)),
			258 => std_logic_vector(to_unsigned(48, 8)),
			259 => std_logic_vector(to_unsigned(239, 8)),
			260 => std_logic_vector(to_unsigned(223, 8)),
			261 => std_logic_vector(to_unsigned(119, 8)),
			262 => std_logic_vector(to_unsigned(227, 8)),
			263 => std_logic_vector(to_unsigned(31, 8)),
			264 => std_logic_vector(to_unsigned(198, 8)),
			265 => std_logic_vector(to_unsigned(80, 8)),
			266 => std_logic_vector(to_unsigned(116, 8)),
			267 => std_logic_vector(to_unsigned(122, 8)),
			268 => std_logic_vector(to_unsigned(116, 8)),
			269 => std_logic_vector(to_unsigned(126, 8)),
			270 => std_logic_vector(to_unsigned(37, 8)),
			271 => std_logic_vector(to_unsigned(210, 8)),
			272 => std_logic_vector(to_unsigned(132, 8)),
			273 => std_logic_vector(to_unsigned(86, 8)),
			274 => std_logic_vector(to_unsigned(123, 8)),
			275 => std_logic_vector(to_unsigned(245, 8)),
			276 => std_logic_vector(to_unsigned(88, 8)),
			277 => std_logic_vector(to_unsigned(183, 8)),
			278 => std_logic_vector(to_unsigned(49, 8)),
			279 => std_logic_vector(to_unsigned(21, 8)),
			280 => std_logic_vector(to_unsigned(146, 8)),
			281 => std_logic_vector(to_unsigned(106, 8)),
			282 => std_logic_vector(to_unsigned(245, 8)),
			283 => std_logic_vector(to_unsigned(214, 8)),
			284 => std_logic_vector(to_unsigned(58, 8)),
			285 => std_logic_vector(to_unsigned(161, 8)),
			286 => std_logic_vector(to_unsigned(221, 8)),
			287 => std_logic_vector(to_unsigned(23, 8)),
			288 => std_logic_vector(to_unsigned(202, 8)),
			289 => std_logic_vector(to_unsigned(98, 8)),
			290 => std_logic_vector(to_unsigned(208, 8)),
			291 => std_logic_vector(to_unsigned(52, 8)),
			292 => std_logic_vector(to_unsigned(141, 8)),
			293 => std_logic_vector(to_unsigned(68, 8)),
			294 => std_logic_vector(to_unsigned(117, 8)),
			295 => std_logic_vector(to_unsigned(244, 8)),
			296 => std_logic_vector(to_unsigned(8, 8)),
			297 => std_logic_vector(to_unsigned(134, 8)),
			298 => std_logic_vector(to_unsigned(10, 8)),
			299 => std_logic_vector(to_unsigned(84, 8)),
			300 => std_logic_vector(to_unsigned(113, 8)),
			301 => std_logic_vector(to_unsigned(43, 8)),
			302 => std_logic_vector(to_unsigned(96, 8)),
			303 => std_logic_vector(to_unsigned(164, 8)),
			304 => std_logic_vector(to_unsigned(34, 8)),
			305 => std_logic_vector(to_unsigned(206, 8)),
			306 => std_logic_vector(to_unsigned(147, 8)),
			307 => std_logic_vector(to_unsigned(6, 8)),
			308 => std_logic_vector(to_unsigned(216, 8)),
			309 => std_logic_vector(to_unsigned(160, 8)),
			310 => std_logic_vector(to_unsigned(115, 8)),
			311 => std_logic_vector(to_unsigned(218, 8)),
			312 => std_logic_vector(to_unsigned(87, 8)),
			313 => std_logic_vector(to_unsigned(249, 8)),
			314 => std_logic_vector(to_unsigned(69, 8)),
			315 => std_logic_vector(to_unsigned(114, 8)),
			316 => std_logic_vector(to_unsigned(164, 8)),
			317 => std_logic_vector(to_unsigned(235, 8)),
			318 => std_logic_vector(to_unsigned(10, 8)),
			319 => std_logic_vector(to_unsigned(245, 8)),
			320 => std_logic_vector(to_unsigned(205, 8)),
			321 => std_logic_vector(to_unsigned(81, 8)),
			322 => std_logic_vector(to_unsigned(22, 8)),
			323 => std_logic_vector(to_unsigned(102, 8)),
			324 => std_logic_vector(to_unsigned(63, 8)),
			325 => std_logic_vector(to_unsigned(33, 8)),
			326 => std_logic_vector(to_unsigned(21, 8)),
			327 => std_logic_vector(to_unsigned(69, 8)),
			328 => std_logic_vector(to_unsigned(185, 8)),
			329 => std_logic_vector(to_unsigned(176, 8)),
			330 => std_logic_vector(to_unsigned(121, 8)),
			331 => std_logic_vector(to_unsigned(121, 8)),
			332 => std_logic_vector(to_unsigned(37, 8)),
			333 => std_logic_vector(to_unsigned(195, 8)),
			334 => std_logic_vector(to_unsigned(25, 8)),
			335 => std_logic_vector(to_unsigned(62, 8)),
			336 => std_logic_vector(to_unsigned(196, 8)),
			337 => std_logic_vector(to_unsigned(91, 8)),
			338 => std_logic_vector(to_unsigned(83, 8)),
			339 => std_logic_vector(to_unsigned(171, 8)),
			340 => std_logic_vector(to_unsigned(29, 8)),
			341 => std_logic_vector(to_unsigned(107, 8)),
			342 => std_logic_vector(to_unsigned(209, 8)),
			343 => std_logic_vector(to_unsigned(174, 8)),
			344 => std_logic_vector(to_unsigned(237, 8)),
			345 => std_logic_vector(to_unsigned(12, 8)),
			346 => std_logic_vector(to_unsigned(121, 8)),
			347 => std_logic_vector(to_unsigned(254, 8)),
			348 => std_logic_vector(to_unsigned(115, 8)),
			349 => std_logic_vector(to_unsigned(2, 8)),
			350 => std_logic_vector(to_unsigned(135, 8)),
			351 => std_logic_vector(to_unsigned(242, 8)),
			352 => std_logic_vector(to_unsigned(101, 8)),
			353 => std_logic_vector(to_unsigned(164, 8)),
			354 => std_logic_vector(to_unsigned(14, 8)),
			355 => std_logic_vector(to_unsigned(105, 8)),
			356 => std_logic_vector(to_unsigned(158, 8)),
			357 => std_logic_vector(to_unsigned(236, 8)),
			358 => std_logic_vector(to_unsigned(184, 8)),
			359 => std_logic_vector(to_unsigned(28, 8)),
			360 => std_logic_vector(to_unsigned(129, 8)),
			361 => std_logic_vector(to_unsigned(27, 8)),
			362 => std_logic_vector(to_unsigned(239, 8)),
			363 => std_logic_vector(to_unsigned(218, 8)),
			364 => std_logic_vector(to_unsigned(188, 8)),
			365 => std_logic_vector(to_unsigned(145, 8)),
			366 => std_logic_vector(to_unsigned(118, 8)),
			367 => std_logic_vector(to_unsigned(112, 8)),
			368 => std_logic_vector(to_unsigned(86, 8)),
			369 => std_logic_vector(to_unsigned(66, 8)),
			370 => std_logic_vector(to_unsigned(214, 8)),
			371 => std_logic_vector(to_unsigned(237, 8)),
			372 => std_logic_vector(to_unsigned(15, 8)),
			373 => std_logic_vector(to_unsigned(152, 8)),
			374 => std_logic_vector(to_unsigned(210, 8)),
			375 => std_logic_vector(to_unsigned(246, 8)),
			376 => std_logic_vector(to_unsigned(165, 8)),
			377 => std_logic_vector(to_unsigned(130, 8)),
			378 => std_logic_vector(to_unsigned(215, 8)),
			379 => std_logic_vector(to_unsigned(118, 8)),
			380 => std_logic_vector(to_unsigned(130, 8)),
			381 => std_logic_vector(to_unsigned(192, 8)),
			382 => std_logic_vector(to_unsigned(40, 8)),
			383 => std_logic_vector(to_unsigned(178, 8)),
			384 => std_logic_vector(to_unsigned(204, 8)),
			385 => std_logic_vector(to_unsigned(101, 8)),
			386 => std_logic_vector(to_unsigned(239, 8)),
			387 => std_logic_vector(to_unsigned(41, 8)),
			388 => std_logic_vector(to_unsigned(188, 8)),
			389 => std_logic_vector(to_unsigned(56, 8)),
			390 => std_logic_vector(to_unsigned(189, 8)),
			391 => std_logic_vector(to_unsigned(134, 8)),
			392 => std_logic_vector(to_unsigned(106, 8)),
			393 => std_logic_vector(to_unsigned(83, 8)),
			394 => std_logic_vector(to_unsigned(253, 8)),
			395 => std_logic_vector(to_unsigned(234, 8)),
			396 => std_logic_vector(to_unsigned(184, 8)),
			397 => std_logic_vector(to_unsigned(90, 8)),
			398 => std_logic_vector(to_unsigned(77, 8)),
			399 => std_logic_vector(to_unsigned(155, 8)),
			400 => std_logic_vector(to_unsigned(162, 8)),
			401 => std_logic_vector(to_unsigned(123, 8)),
			402 => std_logic_vector(to_unsigned(200, 8)),
			403 => std_logic_vector(to_unsigned(151, 8)),
			404 => std_logic_vector(to_unsigned(96, 8)),
			405 => std_logic_vector(to_unsigned(150, 8)),
			406 => std_logic_vector(to_unsigned(28, 8)),
			407 => std_logic_vector(to_unsigned(71, 8)),
			408 => std_logic_vector(to_unsigned(110, 8)),
			409 => std_logic_vector(to_unsigned(44, 8)),
			410 => std_logic_vector(to_unsigned(71, 8)),
			411 => std_logic_vector(to_unsigned(218, 8)),
			412 => std_logic_vector(to_unsigned(167, 8)),
			413 => std_logic_vector(to_unsigned(129, 8)),
			414 => std_logic_vector(to_unsigned(99, 8)),
			415 => std_logic_vector(to_unsigned(225, 8)),
			416 => std_logic_vector(to_unsigned(131, 8)),
			417 => std_logic_vector(to_unsigned(206, 8)),
			418 => std_logic_vector(to_unsigned(143, 8)),
			419 => std_logic_vector(to_unsigned(98, 8)),
			420 => std_logic_vector(to_unsigned(225, 8)),
			421 => std_logic_vector(to_unsigned(127, 8)),
			422 => std_logic_vector(to_unsigned(21, 8)),
			423 => std_logic_vector(to_unsigned(225, 8)),
			424 => std_logic_vector(to_unsigned(149, 8)),
			425 => std_logic_vector(to_unsigned(108, 8)),
			426 => std_logic_vector(to_unsigned(134, 8)),
			427 => std_logic_vector(to_unsigned(90, 8)),
			428 => std_logic_vector(to_unsigned(11, 8)),
			429 => std_logic_vector(to_unsigned(185, 8)),
			430 => std_logic_vector(to_unsigned(106, 8)),
			431 => std_logic_vector(to_unsigned(51, 8)),
			432 => std_logic_vector(to_unsigned(47, 8)),
			433 => std_logic_vector(to_unsigned(229, 8)),
			434 => std_logic_vector(to_unsigned(103, 8)),
			435 => std_logic_vector(to_unsigned(59, 8)),
			436 => std_logic_vector(to_unsigned(6, 8)),
			437 => std_logic_vector(to_unsigned(236, 8)),
			438 => std_logic_vector(to_unsigned(138, 8)),
			439 => std_logic_vector(to_unsigned(28, 8)),
			440 => std_logic_vector(to_unsigned(114, 8)),
			441 => std_logic_vector(to_unsigned(22, 8)),
			442 => std_logic_vector(to_unsigned(209, 8)),
			443 => std_logic_vector(to_unsigned(108, 8)),
			444 => std_logic_vector(to_unsigned(199, 8)),
			445 => std_logic_vector(to_unsigned(215, 8)),
			446 => std_logic_vector(to_unsigned(203, 8)),
			447 => std_logic_vector(to_unsigned(30, 8)),
			448 => std_logic_vector(to_unsigned(246, 8)),
			449 => std_logic_vector(to_unsigned(27, 8)),
			450 => std_logic_vector(to_unsigned(182, 8)),
			451 => std_logic_vector(to_unsigned(132, 8)),
			452 => std_logic_vector(to_unsigned(25, 8)),
			453 => std_logic_vector(to_unsigned(145, 8)),
			454 => std_logic_vector(to_unsigned(174, 8)),
			455 => std_logic_vector(to_unsigned(52, 8)),
			456 => std_logic_vector(to_unsigned(248, 8)),
			457 => std_logic_vector(to_unsigned(196, 8)),
			458 => std_logic_vector(to_unsigned(129, 8)),
			459 => std_logic_vector(to_unsigned(27, 8)),
			460 => std_logic_vector(to_unsigned(46, 8)),
			461 => std_logic_vector(to_unsigned(228, 8)),
			462 => std_logic_vector(to_unsigned(53, 8)),
			463 => std_logic_vector(to_unsigned(136, 8)),
			464 => std_logic_vector(to_unsigned(95, 8)),
			465 => std_logic_vector(to_unsigned(67, 8)),
			466 => std_logic_vector(to_unsigned(228, 8)),
			467 => std_logic_vector(to_unsigned(199, 8)),
			468 => std_logic_vector(to_unsigned(166, 8)),
			469 => std_logic_vector(to_unsigned(138, 8)),
			470 => std_logic_vector(to_unsigned(55, 8)),
			471 => std_logic_vector(to_unsigned(16, 8)),
			472 => std_logic_vector(to_unsigned(22, 8)),
			473 => std_logic_vector(to_unsigned(19, 8)),
			474 => std_logic_vector(to_unsigned(148, 8)),
			475 => std_logic_vector(to_unsigned(187, 8)),
			476 => std_logic_vector(to_unsigned(211, 8)),
			477 => std_logic_vector(to_unsigned(210, 8)),
			478 => std_logic_vector(to_unsigned(81, 8)),
			479 => std_logic_vector(to_unsigned(106, 8)),
			480 => std_logic_vector(to_unsigned(197, 8)),
			481 => std_logic_vector(to_unsigned(243, 8)),
			482 => std_logic_vector(to_unsigned(17, 8)),
			483 => std_logic_vector(to_unsigned(216, 8)),
			484 => std_logic_vector(to_unsigned(233, 8)),
			485 => std_logic_vector(to_unsigned(130, 8)),
			486 => std_logic_vector(to_unsigned(246, 8)),
			487 => std_logic_vector(to_unsigned(80, 8)),
			488 => std_logic_vector(to_unsigned(177, 8)),
			489 => std_logic_vector(to_unsigned(223, 8)),
			490 => std_logic_vector(to_unsigned(193, 8)),
			491 => std_logic_vector(to_unsigned(81, 8)),
			492 => std_logic_vector(to_unsigned(124, 8)),
			493 => std_logic_vector(to_unsigned(6, 8)),
			494 => std_logic_vector(to_unsigned(238, 8)),
			495 => std_logic_vector(to_unsigned(146, 8)),
			496 => std_logic_vector(to_unsigned(163, 8)),
			497 => std_logic_vector(to_unsigned(4, 8)),
			498 => std_logic_vector(to_unsigned(14, 8)),
			499 => std_logic_vector(to_unsigned(27, 8)),
			500 => std_logic_vector(to_unsigned(0, 8)),
			501 => std_logic_vector(to_unsigned(102, 8)),
			502 => std_logic_vector(to_unsigned(197, 8)),
			503 => std_logic_vector(to_unsigned(181, 8)),
			504 => std_logic_vector(to_unsigned(102, 8)),
			505 => std_logic_vector(to_unsigned(114, 8)),
			506 => std_logic_vector(to_unsigned(229, 8)),
			507 => std_logic_vector(to_unsigned(89, 8)),
			508 => std_logic_vector(to_unsigned(102, 8)),
			509 => std_logic_vector(to_unsigned(78, 8)),
			510 => std_logic_vector(to_unsigned(116, 8)),
			511 => std_logic_vector(to_unsigned(248, 8)),
			512 => std_logic_vector(to_unsigned(89, 8)),
			513 => std_logic_vector(to_unsigned(182, 8)),
			514 => std_logic_vector(to_unsigned(64, 8)),
			515 => std_logic_vector(to_unsigned(34, 8)),
			516 => std_logic_vector(to_unsigned(159, 8)),
			517 => std_logic_vector(to_unsigned(209, 8)),
			518 => std_logic_vector(to_unsigned(253, 8)),
			519 => std_logic_vector(to_unsigned(60, 8)),
			520 => std_logic_vector(to_unsigned(98, 8)),
			521 => std_logic_vector(to_unsigned(100, 8)),
			522 => std_logic_vector(to_unsigned(88, 8)),
			523 => std_logic_vector(to_unsigned(250, 8)),
			524 => std_logic_vector(to_unsigned(145, 8)),
			525 => std_logic_vector(to_unsigned(66, 8)),
			526 => std_logic_vector(to_unsigned(197, 8)),
			527 => std_logic_vector(to_unsigned(67, 8)),
			528 => std_logic_vector(to_unsigned(122, 8)),
			529 => std_logic_vector(to_unsigned(62, 8)),
			530 => std_logic_vector(to_unsigned(59, 8)),
			531 => std_logic_vector(to_unsigned(124, 8)),
			532 => std_logic_vector(to_unsigned(36, 8)),
			533 => std_logic_vector(to_unsigned(23, 8)),
			534 => std_logic_vector(to_unsigned(96, 8)),
			535 => std_logic_vector(to_unsigned(131, 8)),
			536 => std_logic_vector(to_unsigned(160, 8)),
			537 => std_logic_vector(to_unsigned(207, 8)),
			538 => std_logic_vector(to_unsigned(92, 8)),
			539 => std_logic_vector(to_unsigned(59, 8)),
			540 => std_logic_vector(to_unsigned(4, 8)),
			541 => std_logic_vector(to_unsigned(248, 8)),
			542 => std_logic_vector(to_unsigned(21, 8)),
			543 => std_logic_vector(to_unsigned(248, 8)),
			544 => std_logic_vector(to_unsigned(91, 8)),
			545 => std_logic_vector(to_unsigned(182, 8)),
			546 => std_logic_vector(to_unsigned(236, 8)),
			547 => std_logic_vector(to_unsigned(139, 8)),
			548 => std_logic_vector(to_unsigned(222, 8)),
			549 => std_logic_vector(to_unsigned(11, 8)),
			550 => std_logic_vector(to_unsigned(99, 8)),
			551 => std_logic_vector(to_unsigned(115, 8)),
			552 => std_logic_vector(to_unsigned(94, 8)),
			553 => std_logic_vector(to_unsigned(17, 8)),
			554 => std_logic_vector(to_unsigned(21, 8)),
			555 => std_logic_vector(to_unsigned(65, 8)),
			556 => std_logic_vector(to_unsigned(206, 8)),
			557 => std_logic_vector(to_unsigned(38, 8)),
			558 => std_logic_vector(to_unsigned(109, 8)),
			559 => std_logic_vector(to_unsigned(62, 8)),
			560 => std_logic_vector(to_unsigned(108, 8)),
			561 => std_logic_vector(to_unsigned(161, 8)),
			562 => std_logic_vector(to_unsigned(46, 8)),
			563 => std_logic_vector(to_unsigned(57, 8)),
			564 => std_logic_vector(to_unsigned(65, 8)),
			565 => std_logic_vector(to_unsigned(153, 8)),
			566 => std_logic_vector(to_unsigned(40, 8)),
			567 => std_logic_vector(to_unsigned(211, 8)),
			568 => std_logic_vector(to_unsigned(69, 8)),
			569 => std_logic_vector(to_unsigned(150, 8)),
			570 => std_logic_vector(to_unsigned(138, 8)),
			571 => std_logic_vector(to_unsigned(24, 8)),
			572 => std_logic_vector(to_unsigned(27, 8)),
			573 => std_logic_vector(to_unsigned(53, 8)),
			574 => std_logic_vector(to_unsigned(9, 8)),
			575 => std_logic_vector(to_unsigned(44, 8)),
			576 => std_logic_vector(to_unsigned(100, 8)),
			577 => std_logic_vector(to_unsigned(48, 8)),
			578 => std_logic_vector(to_unsigned(3, 8)),
			579 => std_logic_vector(to_unsigned(220, 8)),
			580 => std_logic_vector(to_unsigned(211, 8)),
			581 => std_logic_vector(to_unsigned(235, 8)),
			582 => std_logic_vector(to_unsigned(77, 8)),
			583 => std_logic_vector(to_unsigned(75, 8)),
			584 => std_logic_vector(to_unsigned(127, 8)),
			585 => std_logic_vector(to_unsigned(168, 8)),
			586 => std_logic_vector(to_unsigned(129, 8)),
			587 => std_logic_vector(to_unsigned(99, 8)),
			588 => std_logic_vector(to_unsigned(47, 8)),
			589 => std_logic_vector(to_unsigned(105, 8)),
			590 => std_logic_vector(to_unsigned(44, 8)),
			591 => std_logic_vector(to_unsigned(74, 8)),
			592 => std_logic_vector(to_unsigned(6, 8)),
			593 => std_logic_vector(to_unsigned(110, 8)),
			594 => std_logic_vector(to_unsigned(7, 8)),
			595 => std_logic_vector(to_unsigned(30, 8)),
			596 => std_logic_vector(to_unsigned(154, 8)),
			597 => std_logic_vector(to_unsigned(189, 8)),
			598 => std_logic_vector(to_unsigned(56, 8)),
			599 => std_logic_vector(to_unsigned(166, 8)),
			600 => std_logic_vector(to_unsigned(16, 8)),
			601 => std_logic_vector(to_unsigned(147, 8)),
			602 => std_logic_vector(to_unsigned(55, 8)),
			603 => std_logic_vector(to_unsigned(69, 8)),
			604 => std_logic_vector(to_unsigned(225, 8)),
			605 => std_logic_vector(to_unsigned(112, 8)),
			606 => std_logic_vector(to_unsigned(216, 8)),
			607 => std_logic_vector(to_unsigned(249, 8)),
			608 => std_logic_vector(to_unsigned(71, 8)),
			609 => std_logic_vector(to_unsigned(49, 8)),
			610 => std_logic_vector(to_unsigned(160, 8)),
			611 => std_logic_vector(to_unsigned(91, 8)),
			612 => std_logic_vector(to_unsigned(184, 8)),
			613 => std_logic_vector(to_unsigned(25, 8)),
			614 => std_logic_vector(to_unsigned(34, 8)),
			615 => std_logic_vector(to_unsigned(199, 8)),
			616 => std_logic_vector(to_unsigned(92, 8)),
			617 => std_logic_vector(to_unsigned(97, 8)),
			618 => std_logic_vector(to_unsigned(24, 8)),
			619 => std_logic_vector(to_unsigned(120, 8)),
			620 => std_logic_vector(to_unsigned(245, 8)),
			621 => std_logic_vector(to_unsigned(111, 8)),
			622 => std_logic_vector(to_unsigned(58, 8)),
			623 => std_logic_vector(to_unsigned(145, 8)),
			624 => std_logic_vector(to_unsigned(27, 8)),
			625 => std_logic_vector(to_unsigned(59, 8)),
			626 => std_logic_vector(to_unsigned(254, 8)),
			627 => std_logic_vector(to_unsigned(72, 8)),
			628 => std_logic_vector(to_unsigned(29, 8)),
			629 => std_logic_vector(to_unsigned(247, 8)),
			630 => std_logic_vector(to_unsigned(226, 8)),
			631 => std_logic_vector(to_unsigned(175, 8)),
			632 => std_logic_vector(to_unsigned(167, 8)),
			633 => std_logic_vector(to_unsigned(213, 8)),
			634 => std_logic_vector(to_unsigned(97, 8)),
			635 => std_logic_vector(to_unsigned(90, 8)),
			636 => std_logic_vector(to_unsigned(151, 8)),
			637 => std_logic_vector(to_unsigned(28, 8)),
			638 => std_logic_vector(to_unsigned(198, 8)),
			639 => std_logic_vector(to_unsigned(176, 8)),
			640 => std_logic_vector(to_unsigned(73, 8)),
			641 => std_logic_vector(to_unsigned(180, 8)),
			642 => std_logic_vector(to_unsigned(255, 8)),
			643 => std_logic_vector(to_unsigned(192, 8)),
			644 => std_logic_vector(to_unsigned(10, 8)),
			645 => std_logic_vector(to_unsigned(109, 8)),
			646 => std_logic_vector(to_unsigned(14, 8)),
			647 => std_logic_vector(to_unsigned(249, 8)),
			648 => std_logic_vector(to_unsigned(251, 8)),
			649 => std_logic_vector(to_unsigned(72, 8)),
			650 => std_logic_vector(to_unsigned(153, 8)),
			651 => std_logic_vector(to_unsigned(179, 8)),
			652 => std_logic_vector(to_unsigned(101, 8)),
			653 => std_logic_vector(to_unsigned(138, 8)),
			654 => std_logic_vector(to_unsigned(18, 8)),
			655 => std_logic_vector(to_unsigned(82, 8)),
			656 => std_logic_vector(to_unsigned(103, 8)),
			657 => std_logic_vector(to_unsigned(171, 8)),
			658 => std_logic_vector(to_unsigned(13, 8)),
			659 => std_logic_vector(to_unsigned(31, 8)),
			660 => std_logic_vector(to_unsigned(71, 8)),
			661 => std_logic_vector(to_unsigned(128, 8)),
			662 => std_logic_vector(to_unsigned(161, 8)),
			663 => std_logic_vector(to_unsigned(7, 8)),
			664 => std_logic_vector(to_unsigned(104, 8)),
			665 => std_logic_vector(to_unsigned(150, 8)),
			666 => std_logic_vector(to_unsigned(224, 8)),
			667 => std_logic_vector(to_unsigned(159, 8)),
			668 => std_logic_vector(to_unsigned(3, 8)),
			669 => std_logic_vector(to_unsigned(77, 8)),
			670 => std_logic_vector(to_unsigned(239, 8)),
			671 => std_logic_vector(to_unsigned(227, 8)),
			672 => std_logic_vector(to_unsigned(165, 8)),
			673 => std_logic_vector(to_unsigned(106, 8)),
			674 => std_logic_vector(to_unsigned(240, 8)),
			675 => std_logic_vector(to_unsigned(214, 8)),
			676 => std_logic_vector(to_unsigned(90, 8)),
			677 => std_logic_vector(to_unsigned(146, 8)),
			678 => std_logic_vector(to_unsigned(230, 8)),
			679 => std_logic_vector(to_unsigned(245, 8)),
			680 => std_logic_vector(to_unsigned(151, 8)),
			681 => std_logic_vector(to_unsigned(62, 8)),
			682 => std_logic_vector(to_unsigned(23, 8)),
			683 => std_logic_vector(to_unsigned(199, 8)),
			684 => std_logic_vector(to_unsigned(90, 8)),
			685 => std_logic_vector(to_unsigned(210, 8)),
			686 => std_logic_vector(to_unsigned(184, 8)),
			687 => std_logic_vector(to_unsigned(199, 8)),
			688 => std_logic_vector(to_unsigned(163, 8)),
			689 => std_logic_vector(to_unsigned(64, 8)),
			690 => std_logic_vector(to_unsigned(1, 8)),
			691 => std_logic_vector(to_unsigned(4, 8)),
			692 => std_logic_vector(to_unsigned(43, 8)),
			693 => std_logic_vector(to_unsigned(110, 8)),
			694 => std_logic_vector(to_unsigned(211, 8)),
			695 => std_logic_vector(to_unsigned(51, 8)),
			696 => std_logic_vector(to_unsigned(221, 8)),
			697 => std_logic_vector(to_unsigned(211, 8)),
			698 => std_logic_vector(to_unsigned(243, 8)),
			699 => std_logic_vector(to_unsigned(95, 8)),
			700 => std_logic_vector(to_unsigned(132, 8)),
			701 => std_logic_vector(to_unsigned(199, 8)),
			702 => std_logic_vector(to_unsigned(47, 8)),
			703 => std_logic_vector(to_unsigned(197, 8)),
			704 => std_logic_vector(to_unsigned(205, 8)),
			705 => std_logic_vector(to_unsigned(102, 8)),
			706 => std_logic_vector(to_unsigned(178, 8)),
			707 => std_logic_vector(to_unsigned(135, 8)),
			708 => std_logic_vector(to_unsigned(192, 8)),
			709 => std_logic_vector(to_unsigned(34, 8)),
			710 => std_logic_vector(to_unsigned(23, 8)),
			711 => std_logic_vector(to_unsigned(47, 8)),
			712 => std_logic_vector(to_unsigned(66, 8)),
			713 => std_logic_vector(to_unsigned(240, 8)),
			714 => std_logic_vector(to_unsigned(49, 8)),
			715 => std_logic_vector(to_unsigned(42, 8)),
			716 => std_logic_vector(to_unsigned(113, 8)),
			717 => std_logic_vector(to_unsigned(73, 8)),
			718 => std_logic_vector(to_unsigned(58, 8)),
			719 => std_logic_vector(to_unsigned(50, 8)),
			720 => std_logic_vector(to_unsigned(21, 8)),
			721 => std_logic_vector(to_unsigned(9, 8)),
			722 => std_logic_vector(to_unsigned(65, 8)),
			723 => std_logic_vector(to_unsigned(38, 8)),
			724 => std_logic_vector(to_unsigned(161, 8)),
			725 => std_logic_vector(to_unsigned(86, 8)),
			726 => std_logic_vector(to_unsigned(253, 8)),
			727 => std_logic_vector(to_unsigned(12, 8)),
			728 => std_logic_vector(to_unsigned(46, 8)),
			729 => std_logic_vector(to_unsigned(101, 8)),
			730 => std_logic_vector(to_unsigned(16, 8)),
			731 => std_logic_vector(to_unsigned(255, 8)),
			732 => std_logic_vector(to_unsigned(224, 8)),
			733 => std_logic_vector(to_unsigned(181, 8)),
			734 => std_logic_vector(to_unsigned(96, 8)),
			735 => std_logic_vector(to_unsigned(203, 8)),
			736 => std_logic_vector(to_unsigned(134, 8)),
			737 => std_logic_vector(to_unsigned(99, 8)),
			738 => std_logic_vector(to_unsigned(29, 8)),
			739 => std_logic_vector(to_unsigned(216, 8)),
			740 => std_logic_vector(to_unsigned(222, 8)),
			741 => std_logic_vector(to_unsigned(13, 8)),
			742 => std_logic_vector(to_unsigned(156, 8)),
			743 => std_logic_vector(to_unsigned(44, 8)),
			744 => std_logic_vector(to_unsigned(156, 8)),
			745 => std_logic_vector(to_unsigned(70, 8)),
			746 => std_logic_vector(to_unsigned(197, 8)),
			747 => std_logic_vector(to_unsigned(59, 8)),
			748 => std_logic_vector(to_unsigned(58, 8)),
			749 => std_logic_vector(to_unsigned(196, 8)),
			750 => std_logic_vector(to_unsigned(47, 8)),
			751 => std_logic_vector(to_unsigned(201, 8)),
			752 => std_logic_vector(to_unsigned(103, 8)),
			753 => std_logic_vector(to_unsigned(27, 8)),
			754 => std_logic_vector(to_unsigned(146, 8)),
			755 => std_logic_vector(to_unsigned(237, 8)),
			756 => std_logic_vector(to_unsigned(58, 8)),
			757 => std_logic_vector(to_unsigned(60, 8)),
			758 => std_logic_vector(to_unsigned(85, 8)),
			759 => std_logic_vector(to_unsigned(158, 8)),
			760 => std_logic_vector(to_unsigned(142, 8)),
			761 => std_logic_vector(to_unsigned(95, 8)),
			762 => std_logic_vector(to_unsigned(52, 8)),
			763 => std_logic_vector(to_unsigned(64, 8)),
			764 => std_logic_vector(to_unsigned(41, 8)),
			765 => std_logic_vector(to_unsigned(95, 8)),
			766 => std_logic_vector(to_unsigned(145, 8)),
			767 => std_logic_vector(to_unsigned(173, 8)),
			768 => std_logic_vector(to_unsigned(35, 8)),
			769 => std_logic_vector(to_unsigned(14, 8)),
			770 => std_logic_vector(to_unsigned(231, 8)),
			771 => std_logic_vector(to_unsigned(70, 8)),
			772 => std_logic_vector(to_unsigned(184, 8)),
			773 => std_logic_vector(to_unsigned(192, 8)),
			774 => std_logic_vector(to_unsigned(207, 8)),
			775 => std_logic_vector(to_unsigned(153, 8)),
			776 => std_logic_vector(to_unsigned(185, 8)),
			777 => std_logic_vector(to_unsigned(134, 8)),
			778 => std_logic_vector(to_unsigned(239, 8)),
			779 => std_logic_vector(to_unsigned(241, 8)),
			780 => std_logic_vector(to_unsigned(230, 8)),
			781 => std_logic_vector(to_unsigned(234, 8)),
			782 => std_logic_vector(to_unsigned(19, 8)),
			783 => std_logic_vector(to_unsigned(144, 8)),
			784 => std_logic_vector(to_unsigned(68, 8)),
			785 => std_logic_vector(to_unsigned(8, 8)),
			786 => std_logic_vector(to_unsigned(115, 8)),
			787 => std_logic_vector(to_unsigned(30, 8)),
			788 => std_logic_vector(to_unsigned(172, 8)),
			789 => std_logic_vector(to_unsigned(42, 8)),
			790 => std_logic_vector(to_unsigned(129, 8)),
			791 => std_logic_vector(to_unsigned(172, 8)),
			792 => std_logic_vector(to_unsigned(69, 8)),
			793 => std_logic_vector(to_unsigned(136, 8)),
			794 => std_logic_vector(to_unsigned(206, 8)),
			795 => std_logic_vector(to_unsigned(139, 8)),
			796 => std_logic_vector(to_unsigned(77, 8)),
			797 => std_logic_vector(to_unsigned(142, 8)),
			798 => std_logic_vector(to_unsigned(153, 8)),
			799 => std_logic_vector(to_unsigned(198, 8)),
			800 => std_logic_vector(to_unsigned(24, 8)),
			801 => std_logic_vector(to_unsigned(225, 8)),
			802 => std_logic_vector(to_unsigned(132, 8)),
			803 => std_logic_vector(to_unsigned(9, 8)),
			804 => std_logic_vector(to_unsigned(50, 8)),
			805 => std_logic_vector(to_unsigned(209, 8)),
			806 => std_logic_vector(to_unsigned(111, 8)),
			807 => std_logic_vector(to_unsigned(120, 8)),
			808 => std_logic_vector(to_unsigned(32, 8)),
			809 => std_logic_vector(to_unsigned(4, 8)),
			810 => std_logic_vector(to_unsigned(39, 8)),
			811 => std_logic_vector(to_unsigned(237, 8)),
			812 => std_logic_vector(to_unsigned(183, 8)),
			813 => std_logic_vector(to_unsigned(94, 8)),
			814 => std_logic_vector(to_unsigned(220, 8)),
			815 => std_logic_vector(to_unsigned(104, 8)),
			816 => std_logic_vector(to_unsigned(190, 8)),
			817 => std_logic_vector(to_unsigned(40, 8)),
			818 => std_logic_vector(to_unsigned(105, 8)),
			819 => std_logic_vector(to_unsigned(189, 8)),
			820 => std_logic_vector(to_unsigned(98, 8)),
			821 => std_logic_vector(to_unsigned(186, 8)),
			822 => std_logic_vector(to_unsigned(221, 8)),
			823 => std_logic_vector(to_unsigned(194, 8)),
			824 => std_logic_vector(to_unsigned(237, 8)),
			825 => std_logic_vector(to_unsigned(7, 8)),
			826 => std_logic_vector(to_unsigned(33, 8)),
			827 => std_logic_vector(to_unsigned(134, 8)),
			828 => std_logic_vector(to_unsigned(162, 8)),
			829 => std_logic_vector(to_unsigned(152, 8)),
			830 => std_logic_vector(to_unsigned(203, 8)),
			831 => std_logic_vector(to_unsigned(232, 8)),
			832 => std_logic_vector(to_unsigned(207, 8)),
			833 => std_logic_vector(to_unsigned(74, 8)),
			834 => std_logic_vector(to_unsigned(147, 8)),
			835 => std_logic_vector(to_unsigned(183, 8)),
			836 => std_logic_vector(to_unsigned(69, 8)),
			837 => std_logic_vector(to_unsigned(27, 8)),
			838 => std_logic_vector(to_unsigned(94, 8)),
			839 => std_logic_vector(to_unsigned(34, 8)),
			840 => std_logic_vector(to_unsigned(135, 8)),
			841 => std_logic_vector(to_unsigned(148, 8)),
			842 => std_logic_vector(to_unsigned(45, 8)),
			843 => std_logic_vector(to_unsigned(187, 8)),
			844 => std_logic_vector(to_unsigned(241, 8)),
			845 => std_logic_vector(to_unsigned(160, 8)),
			846 => std_logic_vector(to_unsigned(177, 8)),
			847 => std_logic_vector(to_unsigned(30, 8)),
			848 => std_logic_vector(to_unsigned(206, 8)),
			849 => std_logic_vector(to_unsigned(113, 8)),
			850 => std_logic_vector(to_unsigned(181, 8)),
			851 => std_logic_vector(to_unsigned(112, 8)),
			852 => std_logic_vector(to_unsigned(159, 8)),
			853 => std_logic_vector(to_unsigned(74, 8)),
			854 => std_logic_vector(to_unsigned(108, 8)),
			855 => std_logic_vector(to_unsigned(185, 8)),
			856 => std_logic_vector(to_unsigned(121, 8)),
			857 => std_logic_vector(to_unsigned(187, 8)),
			858 => std_logic_vector(to_unsigned(42, 8)),
			859 => std_logic_vector(to_unsigned(247, 8)),
			860 => std_logic_vector(to_unsigned(238, 8)),
			861 => std_logic_vector(to_unsigned(112, 8)),
			862 => std_logic_vector(to_unsigned(209, 8)),
			863 => std_logic_vector(to_unsigned(29, 8)),
			864 => std_logic_vector(to_unsigned(251, 8)),
			865 => std_logic_vector(to_unsigned(217, 8)),
			866 => std_logic_vector(to_unsigned(32, 8)),
			867 => std_logic_vector(to_unsigned(206, 8)),
			868 => std_logic_vector(to_unsigned(247, 8)),
			869 => std_logic_vector(to_unsigned(63, 8)),
			870 => std_logic_vector(to_unsigned(212, 8)),
			871 => std_logic_vector(to_unsigned(194, 8)),
			872 => std_logic_vector(to_unsigned(201, 8)),
			873 => std_logic_vector(to_unsigned(230, 8)),
			874 => std_logic_vector(to_unsigned(182, 8)),
			875 => std_logic_vector(to_unsigned(234, 8)),
			876 => std_logic_vector(to_unsigned(42, 8)),
			877 => std_logic_vector(to_unsigned(40, 8)),
			878 => std_logic_vector(to_unsigned(25, 8)),
			879 => std_logic_vector(to_unsigned(120, 8)),
			880 => std_logic_vector(to_unsigned(137, 8)),
			881 => std_logic_vector(to_unsigned(233, 8)),
			882 => std_logic_vector(to_unsigned(75, 8)),
			883 => std_logic_vector(to_unsigned(150, 8)),
			884 => std_logic_vector(to_unsigned(133, 8)),
			885 => std_logic_vector(to_unsigned(223, 8)),
			886 => std_logic_vector(to_unsigned(66, 8)),
			887 => std_logic_vector(to_unsigned(40, 8)),
			888 => std_logic_vector(to_unsigned(237, 8)),
			889 => std_logic_vector(to_unsigned(74, 8)),
			890 => std_logic_vector(to_unsigned(74, 8)),
			891 => std_logic_vector(to_unsigned(150, 8)),
			892 => std_logic_vector(to_unsigned(237, 8)),
			893 => std_logic_vector(to_unsigned(236, 8)),
			894 => std_logic_vector(to_unsigned(218, 8)),
			895 => std_logic_vector(to_unsigned(10, 8)),
			896 => std_logic_vector(to_unsigned(68, 8)),
			897 => std_logic_vector(to_unsigned(181, 8)),
			898 => std_logic_vector(to_unsigned(102, 8)),
			899 => std_logic_vector(to_unsigned(191, 8)),
			900 => std_logic_vector(to_unsigned(173, 8)),
			901 => std_logic_vector(to_unsigned(159, 8)),
			902 => std_logic_vector(to_unsigned(236, 8)),
			903 => std_logic_vector(to_unsigned(157, 8)),
			904 => std_logic_vector(to_unsigned(142, 8)),
			905 => std_logic_vector(to_unsigned(174, 8)),
			906 => std_logic_vector(to_unsigned(130, 8)),
			907 => std_logic_vector(to_unsigned(65, 8)),
			908 => std_logic_vector(to_unsigned(181, 8)),
			909 => std_logic_vector(to_unsigned(193, 8)),
			910 => std_logic_vector(to_unsigned(161, 8)),
			911 => std_logic_vector(to_unsigned(25, 8)),
			912 => std_logic_vector(to_unsigned(220, 8)),
			913 => std_logic_vector(to_unsigned(190, 8)),
			914 => std_logic_vector(to_unsigned(78, 8)),
			915 => std_logic_vector(to_unsigned(109, 8)),
			916 => std_logic_vector(to_unsigned(72, 8)),
			917 => std_logic_vector(to_unsigned(135, 8)),
			918 => std_logic_vector(to_unsigned(106, 8)),
			919 => std_logic_vector(to_unsigned(193, 8)),
			920 => std_logic_vector(to_unsigned(197, 8)),
			921 => std_logic_vector(to_unsigned(59, 8)),
			922 => std_logic_vector(to_unsigned(253, 8)),
			923 => std_logic_vector(to_unsigned(166, 8)),
			924 => std_logic_vector(to_unsigned(23, 8)),
			925 => std_logic_vector(to_unsigned(183, 8)),
			926 => std_logic_vector(to_unsigned(221, 8)),
			927 => std_logic_vector(to_unsigned(164, 8)),
			928 => std_logic_vector(to_unsigned(233, 8)),
			929 => std_logic_vector(to_unsigned(15, 8)),
			930 => std_logic_vector(to_unsigned(15, 8)),
			931 => std_logic_vector(to_unsigned(1, 8)),
			932 => std_logic_vector(to_unsigned(44, 8)),
			933 => std_logic_vector(to_unsigned(58, 8)),
			934 => std_logic_vector(to_unsigned(126, 8)),
			935 => std_logic_vector(to_unsigned(222, 8)),
			936 => std_logic_vector(to_unsigned(167, 8)),
			937 => std_logic_vector(to_unsigned(225, 8)),
			938 => std_logic_vector(to_unsigned(193, 8)),
			939 => std_logic_vector(to_unsigned(215, 8)),
			940 => std_logic_vector(to_unsigned(187, 8)),
			941 => std_logic_vector(to_unsigned(234, 8)),
			942 => std_logic_vector(to_unsigned(221, 8)),
			943 => std_logic_vector(to_unsigned(47, 8)),
			944 => std_logic_vector(to_unsigned(162, 8)),
			945 => std_logic_vector(to_unsigned(7, 8)),
			946 => std_logic_vector(to_unsigned(34, 8)),
			947 => std_logic_vector(to_unsigned(1, 8)),
			948 => std_logic_vector(to_unsigned(167, 8)),
			949 => std_logic_vector(to_unsigned(234, 8)),
			950 => std_logic_vector(to_unsigned(163, 8)),
			951 => std_logic_vector(to_unsigned(195, 8)),
			952 => std_logic_vector(to_unsigned(245, 8)),
			953 => std_logic_vector(to_unsigned(75, 8)),
			954 => std_logic_vector(to_unsigned(191, 8)),
			955 => std_logic_vector(to_unsigned(168, 8)),
			956 => std_logic_vector(to_unsigned(245, 8)),
			957 => std_logic_vector(to_unsigned(191, 8)),
			958 => std_logic_vector(to_unsigned(43, 8)),
			959 => std_logic_vector(to_unsigned(195, 8)),
			960 => std_logic_vector(to_unsigned(150, 8)),
			961 => std_logic_vector(to_unsigned(130, 8)),
			962 => std_logic_vector(to_unsigned(177, 8)),
			963 => std_logic_vector(to_unsigned(130, 8)),
			964 => std_logic_vector(to_unsigned(124, 8)),
			965 => std_logic_vector(to_unsigned(211, 8)),
			966 => std_logic_vector(to_unsigned(190, 8)),
			967 => std_logic_vector(to_unsigned(76, 8)),
			968 => std_logic_vector(to_unsigned(37, 8)),
			969 => std_logic_vector(to_unsigned(5, 8)),
			970 => std_logic_vector(to_unsigned(77, 8)),
			971 => std_logic_vector(to_unsigned(0, 8)),
			972 => std_logic_vector(to_unsigned(215, 8)),
			973 => std_logic_vector(to_unsigned(3, 8)),
			974 => std_logic_vector(to_unsigned(35, 8)),
			975 => std_logic_vector(to_unsigned(219, 8)),
			976 => std_logic_vector(to_unsigned(156, 8)),
			977 => std_logic_vector(to_unsigned(240, 8)),
			978 => std_logic_vector(to_unsigned(90, 8)),
			979 => std_logic_vector(to_unsigned(15, 8)),
			980 => std_logic_vector(to_unsigned(216, 8)),
			981 => std_logic_vector(to_unsigned(47, 8)),
			982 => std_logic_vector(to_unsigned(122, 8)),
			983 => std_logic_vector(to_unsigned(107, 8)),
			984 => std_logic_vector(to_unsigned(85, 8)),
			985 => std_logic_vector(to_unsigned(103, 8)),
			986 => std_logic_vector(to_unsigned(42, 8)),
			987 => std_logic_vector(to_unsigned(15, 8)),
			988 => std_logic_vector(to_unsigned(133, 8)),
			989 => std_logic_vector(to_unsigned(170, 8)),
			990 => std_logic_vector(to_unsigned(143, 8)),
			991 => std_logic_vector(to_unsigned(73, 8)),
			992 => std_logic_vector(to_unsigned(116, 8)),
			993 => std_logic_vector(to_unsigned(137, 8)),
			994 => std_logic_vector(to_unsigned(221, 8)),
			995 => std_logic_vector(to_unsigned(79, 8)),
			996 => std_logic_vector(to_unsigned(254, 8)),
			997 => std_logic_vector(to_unsigned(162, 8)),
			998 => std_logic_vector(to_unsigned(242, 8)),
			999 => std_logic_vector(to_unsigned(87, 8)),
			1000 => std_logic_vector(to_unsigned(3, 8)),
			1001 => std_logic_vector(to_unsigned(222, 8)),
			1002 => std_logic_vector(to_unsigned(97, 8)),
			1003 => std_logic_vector(to_unsigned(170, 8)),
			1004 => std_logic_vector(to_unsigned(71, 8)),
			1005 => std_logic_vector(to_unsigned(223, 8)),
			1006 => std_logic_vector(to_unsigned(13, 8)),
			1007 => std_logic_vector(to_unsigned(229, 8)),
			1008 => std_logic_vector(to_unsigned(140, 8)),
			1009 => std_logic_vector(to_unsigned(193, 8)),
			1010 => std_logic_vector(to_unsigned(238, 8)),
			1011 => std_logic_vector(to_unsigned(54, 8)),
			1012 => std_logic_vector(to_unsigned(220, 8)),
			1013 => std_logic_vector(to_unsigned(86, 8)),
			1014 => std_logic_vector(to_unsigned(235, 8)),
			1015 => std_logic_vector(to_unsigned(202, 8)),
			1016 => std_logic_vector(to_unsigned(93, 8)),
			1017 => std_logic_vector(to_unsigned(73, 8)),
			1018 => std_logic_vector(to_unsigned(78, 8)),
			1019 => std_logic_vector(to_unsigned(43, 8)),
			1020 => std_logic_vector(to_unsigned(185, 8)),
			1021 => std_logic_vector(to_unsigned(163, 8)),
			1022 => std_logic_vector(to_unsigned(244, 8)),
			1023 => std_logic_vector(to_unsigned(130, 8)),
			1024 => std_logic_vector(to_unsigned(145, 8)),
			1025 => std_logic_vector(to_unsigned(235, 8)),
			1026 => std_logic_vector(to_unsigned(61, 8)),
			1027 => std_logic_vector(to_unsigned(77, 8)),
			1028 => std_logic_vector(to_unsigned(225, 8)),
			1029 => std_logic_vector(to_unsigned(125, 8)),
			1030 => std_logic_vector(to_unsigned(35, 8)),
			1031 => std_logic_vector(to_unsigned(228, 8)),
			1032 => std_logic_vector(to_unsigned(250, 8)),
			1033 => std_logic_vector(to_unsigned(41, 8)),
			1034 => std_logic_vector(to_unsigned(215, 8)),
			1035 => std_logic_vector(to_unsigned(253, 8)),
			1036 => std_logic_vector(to_unsigned(58, 8)),
			1037 => std_logic_vector(to_unsigned(128, 8)),
			1038 => std_logic_vector(to_unsigned(98, 8)),
			1039 => std_logic_vector(to_unsigned(24, 8)),
			1040 => std_logic_vector(to_unsigned(191, 8)),
			1041 => std_logic_vector(to_unsigned(216, 8)),
			1042 => std_logic_vector(to_unsigned(127, 8)),
			1043 => std_logic_vector(to_unsigned(44, 8)),
			1044 => std_logic_vector(to_unsigned(91, 8)),
			1045 => std_logic_vector(to_unsigned(9, 8)),
			1046 => std_logic_vector(to_unsigned(42, 8)),
			1047 => std_logic_vector(to_unsigned(208, 8)),
			1048 => std_logic_vector(to_unsigned(239, 8)),
			1049 => std_logic_vector(to_unsigned(187, 8)),
			1050 => std_logic_vector(to_unsigned(213, 8)),
			1051 => std_logic_vector(to_unsigned(117, 8)),
			1052 => std_logic_vector(to_unsigned(211, 8)),
			1053 => std_logic_vector(to_unsigned(158, 8)),
			1054 => std_logic_vector(to_unsigned(191, 8)),
			1055 => std_logic_vector(to_unsigned(62, 8)),
			1056 => std_logic_vector(to_unsigned(254, 8)),
			1057 => std_logic_vector(to_unsigned(117, 8)),
			1058 => std_logic_vector(to_unsigned(86, 8)),
			1059 => std_logic_vector(to_unsigned(245, 8)),
			1060 => std_logic_vector(to_unsigned(167, 8)),
			1061 => std_logic_vector(to_unsigned(169, 8)),
			1062 => std_logic_vector(to_unsigned(51, 8)),
			1063 => std_logic_vector(to_unsigned(217, 8)),
			1064 => std_logic_vector(to_unsigned(233, 8)),
			1065 => std_logic_vector(to_unsigned(254, 8)),
			1066 => std_logic_vector(to_unsigned(120, 8)),
			1067 => std_logic_vector(to_unsigned(19, 8)),
			1068 => std_logic_vector(to_unsigned(213, 8)),
			1069 => std_logic_vector(to_unsigned(125, 8)),
			1070 => std_logic_vector(to_unsigned(239, 8)),
			1071 => std_logic_vector(to_unsigned(147, 8)),
			1072 => std_logic_vector(to_unsigned(206, 8)),
			1073 => std_logic_vector(to_unsigned(19, 8)),
			1074 => std_logic_vector(to_unsigned(255, 8)),
			1075 => std_logic_vector(to_unsigned(172, 8)),
			1076 => std_logic_vector(to_unsigned(49, 8)),
			1077 => std_logic_vector(to_unsigned(217, 8)),
			1078 => std_logic_vector(to_unsigned(147, 8)),
			1079 => std_logic_vector(to_unsigned(97, 8)),
			1080 => std_logic_vector(to_unsigned(30, 8)),
			1081 => std_logic_vector(to_unsigned(80, 8)),
			1082 => std_logic_vector(to_unsigned(37, 8)),
			1083 => std_logic_vector(to_unsigned(143, 8)),
			1084 => std_logic_vector(to_unsigned(31, 8)),
			1085 => std_logic_vector(to_unsigned(129, 8)),
			1086 => std_logic_vector(to_unsigned(13, 8)),
			1087 => std_logic_vector(to_unsigned(118, 8)),
			1088 => std_logic_vector(to_unsigned(169, 8)),
			1089 => std_logic_vector(to_unsigned(249, 8)),
			1090 => std_logic_vector(to_unsigned(225, 8)),
			1091 => std_logic_vector(to_unsigned(97, 8)),
			1092 => std_logic_vector(to_unsigned(17, 8)),
			1093 => std_logic_vector(to_unsigned(100, 8)),
			1094 => std_logic_vector(to_unsigned(70, 8)),
			1095 => std_logic_vector(to_unsigned(64, 8)),
			1096 => std_logic_vector(to_unsigned(0, 8)),
			1097 => std_logic_vector(to_unsigned(208, 8)),
			1098 => std_logic_vector(to_unsigned(240, 8)),
			1099 => std_logic_vector(to_unsigned(20, 8)),
			1100 => std_logic_vector(to_unsigned(245, 8)),
			1101 => std_logic_vector(to_unsigned(123, 8)),
			1102 => std_logic_vector(to_unsigned(170, 8)),
			1103 => std_logic_vector(to_unsigned(141, 8)),
			1104 => std_logic_vector(to_unsigned(1, 8)),
			1105 => std_logic_vector(to_unsigned(231, 8)),
			1106 => std_logic_vector(to_unsigned(102, 8)),
			1107 => std_logic_vector(to_unsigned(255, 8)),
			1108 => std_logic_vector(to_unsigned(32, 8)),
			1109 => std_logic_vector(to_unsigned(16, 8)),
			1110 => std_logic_vector(to_unsigned(254, 8)),
			1111 => std_logic_vector(to_unsigned(121, 8)),
			1112 => std_logic_vector(to_unsigned(194, 8)),
			1113 => std_logic_vector(to_unsigned(149, 8)),
			1114 => std_logic_vector(to_unsigned(117, 8)),
			1115 => std_logic_vector(to_unsigned(51, 8)),
			1116 => std_logic_vector(to_unsigned(41, 8)),
			1117 => std_logic_vector(to_unsigned(90, 8)),
			1118 => std_logic_vector(to_unsigned(228, 8)),
			1119 => std_logic_vector(to_unsigned(107, 8)),
			1120 => std_logic_vector(to_unsigned(111, 8)),
			1121 => std_logic_vector(to_unsigned(44, 8)),
			1122 => std_logic_vector(to_unsigned(113, 8)),
			1123 => std_logic_vector(to_unsigned(138, 8)),
			1124 => std_logic_vector(to_unsigned(109, 8)),
			1125 => std_logic_vector(to_unsigned(177, 8)),
			1126 => std_logic_vector(to_unsigned(238, 8)),
			1127 => std_logic_vector(to_unsigned(188, 8)),
			1128 => std_logic_vector(to_unsigned(107, 8)),
			1129 => std_logic_vector(to_unsigned(219, 8)),
			1130 => std_logic_vector(to_unsigned(41, 8)),
			1131 => std_logic_vector(to_unsigned(193, 8)),
			1132 => std_logic_vector(to_unsigned(153, 8)),
			1133 => std_logic_vector(to_unsigned(249, 8)),
			1134 => std_logic_vector(to_unsigned(79, 8)),
			1135 => std_logic_vector(to_unsigned(225, 8)),
			1136 => std_logic_vector(to_unsigned(71, 8)),
			1137 => std_logic_vector(to_unsigned(34, 8)),
			1138 => std_logic_vector(to_unsigned(196, 8)),
			1139 => std_logic_vector(to_unsigned(183, 8)),
			1140 => std_logic_vector(to_unsigned(168, 8)),
			1141 => std_logic_vector(to_unsigned(212, 8)),
			1142 => std_logic_vector(to_unsigned(48, 8)),
			1143 => std_logic_vector(to_unsigned(135, 8)),
			1144 => std_logic_vector(to_unsigned(22, 8)),
			1145 => std_logic_vector(to_unsigned(100, 8)),
			1146 => std_logic_vector(to_unsigned(208, 8)),
			1147 => std_logic_vector(to_unsigned(230, 8)),
			1148 => std_logic_vector(to_unsigned(78, 8)),
			1149 => std_logic_vector(to_unsigned(72, 8)),
			1150 => std_logic_vector(to_unsigned(172, 8)),
			1151 => std_logic_vector(to_unsigned(203, 8)),
			1152 => std_logic_vector(to_unsigned(189, 8)),
			1153 => std_logic_vector(to_unsigned(197, 8)),
			1154 => std_logic_vector(to_unsigned(241, 8)),
			1155 => std_logic_vector(to_unsigned(129, 8)),
			1156 => std_logic_vector(to_unsigned(84, 8)),
			1157 => std_logic_vector(to_unsigned(162, 8)),
			1158 => std_logic_vector(to_unsigned(36, 8)),
			1159 => std_logic_vector(to_unsigned(255, 8)),
			1160 => std_logic_vector(to_unsigned(169, 8)),
			1161 => std_logic_vector(to_unsigned(36, 8)),
			1162 => std_logic_vector(to_unsigned(248, 8)),
			1163 => std_logic_vector(to_unsigned(162, 8)),
			1164 => std_logic_vector(to_unsigned(10, 8)),
			1165 => std_logic_vector(to_unsigned(152, 8)),
			1166 => std_logic_vector(to_unsigned(41, 8)),
			1167 => std_logic_vector(to_unsigned(89, 8)),
			1168 => std_logic_vector(to_unsigned(104, 8)),
			1169 => std_logic_vector(to_unsigned(49, 8)),
			1170 => std_logic_vector(to_unsigned(175, 8)),
			1171 => std_logic_vector(to_unsigned(64, 8)),
			1172 => std_logic_vector(to_unsigned(51, 8)),
			1173 => std_logic_vector(to_unsigned(129, 8)),
			1174 => std_logic_vector(to_unsigned(124, 8)),
			1175 => std_logic_vector(to_unsigned(15, 8)),
			1176 => std_logic_vector(to_unsigned(25, 8)),
			1177 => std_logic_vector(to_unsigned(82, 8)),
			1178 => std_logic_vector(to_unsigned(149, 8)),
			1179 => std_logic_vector(to_unsigned(184, 8)),
			1180 => std_logic_vector(to_unsigned(38, 8)),
			1181 => std_logic_vector(to_unsigned(232, 8)),
			1182 => std_logic_vector(to_unsigned(87, 8)),
			1183 => std_logic_vector(to_unsigned(211, 8)),
			1184 => std_logic_vector(to_unsigned(166, 8)),
			1185 => std_logic_vector(to_unsigned(33, 8)),
			1186 => std_logic_vector(to_unsigned(5, 8)),
			1187 => std_logic_vector(to_unsigned(156, 8)),
			1188 => std_logic_vector(to_unsigned(3, 8)),
			1189 => std_logic_vector(to_unsigned(173, 8)),
			1190 => std_logic_vector(to_unsigned(100, 8)),
			1191 => std_logic_vector(to_unsigned(59, 8)),
			1192 => std_logic_vector(to_unsigned(88, 8)),
			1193 => std_logic_vector(to_unsigned(67, 8)),
			1194 => std_logic_vector(to_unsigned(205, 8)),
			1195 => std_logic_vector(to_unsigned(161, 8)),
			1196 => std_logic_vector(to_unsigned(112, 8)),
			1197 => std_logic_vector(to_unsigned(105, 8)),
			1198 => std_logic_vector(to_unsigned(176, 8)),
			1199 => std_logic_vector(to_unsigned(131, 8)),
			1200 => std_logic_vector(to_unsigned(119, 8)),
			1201 => std_logic_vector(to_unsigned(59, 8)),
			1202 => std_logic_vector(to_unsigned(105, 8)),
			1203 => std_logic_vector(to_unsigned(237, 8)),
			1204 => std_logic_vector(to_unsigned(83, 8)),
			1205 => std_logic_vector(to_unsigned(145, 8)),
			1206 => std_logic_vector(to_unsigned(253, 8)),
			1207 => std_logic_vector(to_unsigned(50, 8)),
			1208 => std_logic_vector(to_unsigned(179, 8)),
			1209 => std_logic_vector(to_unsigned(66, 8)),
			1210 => std_logic_vector(to_unsigned(153, 8)),
			1211 => std_logic_vector(to_unsigned(137, 8)),
			1212 => std_logic_vector(to_unsigned(158, 8)),
			1213 => std_logic_vector(to_unsigned(239, 8)),
			1214 => std_logic_vector(to_unsigned(121, 8)),
			1215 => std_logic_vector(to_unsigned(82, 8)),
			1216 => std_logic_vector(to_unsigned(128, 8)),
			1217 => std_logic_vector(to_unsigned(208, 8)),
			1218 => std_logic_vector(to_unsigned(156, 8)),
			1219 => std_logic_vector(to_unsigned(66, 8)),
			1220 => std_logic_vector(to_unsigned(181, 8)),
			1221 => std_logic_vector(to_unsigned(115, 8)),
			1222 => std_logic_vector(to_unsigned(44, 8)),
			1223 => std_logic_vector(to_unsigned(111, 8)),
			1224 => std_logic_vector(to_unsigned(232, 8)),
			1225 => std_logic_vector(to_unsigned(190, 8)),
			1226 => std_logic_vector(to_unsigned(212, 8)),
			1227 => std_logic_vector(to_unsigned(127, 8)),
			1228 => std_logic_vector(to_unsigned(147, 8)),
			1229 => std_logic_vector(to_unsigned(212, 8)),
			1230 => std_logic_vector(to_unsigned(131, 8)),
			1231 => std_logic_vector(to_unsigned(214, 8)),
			1232 => std_logic_vector(to_unsigned(195, 8)),
			1233 => std_logic_vector(to_unsigned(37, 8)),
			1234 => std_logic_vector(to_unsigned(250, 8)),
			1235 => std_logic_vector(to_unsigned(86, 8)),
			1236 => std_logic_vector(to_unsigned(180, 8)),
			1237 => std_logic_vector(to_unsigned(189, 8)),
			1238 => std_logic_vector(to_unsigned(188, 8)),
			1239 => std_logic_vector(to_unsigned(85, 8)),
			1240 => std_logic_vector(to_unsigned(228, 8)),
			1241 => std_logic_vector(to_unsigned(67, 8)),
			1242 => std_logic_vector(to_unsigned(178, 8)),
			1243 => std_logic_vector(to_unsigned(19, 8)),
			1244 => std_logic_vector(to_unsigned(200, 8)),
			1245 => std_logic_vector(to_unsigned(120, 8)),
			1246 => std_logic_vector(to_unsigned(9, 8)),
			1247 => std_logic_vector(to_unsigned(42, 8)),
			1248 => std_logic_vector(to_unsigned(250, 8)),
			1249 => std_logic_vector(to_unsigned(215, 8)),
			1250 => std_logic_vector(to_unsigned(18, 8)),
			1251 => std_logic_vector(to_unsigned(139, 8)),
			1252 => std_logic_vector(to_unsigned(14, 8)),
			1253 => std_logic_vector(to_unsigned(202, 8)),
			1254 => std_logic_vector(to_unsigned(36, 8)),
			1255 => std_logic_vector(to_unsigned(140, 8)),
			1256 => std_logic_vector(to_unsigned(115, 8)),
			1257 => std_logic_vector(to_unsigned(254, 8)),
			1258 => std_logic_vector(to_unsigned(89, 8)),
			1259 => std_logic_vector(to_unsigned(149, 8)),
			1260 => std_logic_vector(to_unsigned(32, 8)),
			1261 => std_logic_vector(to_unsigned(47, 8)),
			1262 => std_logic_vector(to_unsigned(102, 8)),
			1263 => std_logic_vector(to_unsigned(164, 8)),
			1264 => std_logic_vector(to_unsigned(249, 8)),
			1265 => std_logic_vector(to_unsigned(58, 8)),
			1266 => std_logic_vector(to_unsigned(151, 8)),
			1267 => std_logic_vector(to_unsigned(112, 8)),
			1268 => std_logic_vector(to_unsigned(134, 8)),
			1269 => std_logic_vector(to_unsigned(99, 8)),
			1270 => std_logic_vector(to_unsigned(2, 8)),
			1271 => std_logic_vector(to_unsigned(8, 8)),
			1272 => std_logic_vector(to_unsigned(246, 8)),
			1273 => std_logic_vector(to_unsigned(208, 8)),
			1274 => std_logic_vector(to_unsigned(216, 8)),
			1275 => std_logic_vector(to_unsigned(89, 8)),
			1276 => std_logic_vector(to_unsigned(191, 8)),
			1277 => std_logic_vector(to_unsigned(109, 8)),
			1278 => std_logic_vector(to_unsigned(163, 8)),
			1279 => std_logic_vector(to_unsigned(76, 8)),
			1280 => std_logic_vector(to_unsigned(63, 8)),
			1281 => std_logic_vector(to_unsigned(56, 8)),
			1282 => std_logic_vector(to_unsigned(7, 8)),
			1283 => std_logic_vector(to_unsigned(17, 8)),
			1284 => std_logic_vector(to_unsigned(218, 8)),
			1285 => std_logic_vector(to_unsigned(223, 8)),
			1286 => std_logic_vector(to_unsigned(164, 8)),
			1287 => std_logic_vector(to_unsigned(162, 8)),
			1288 => std_logic_vector(to_unsigned(110, 8)),
			1289 => std_logic_vector(to_unsigned(229, 8)),
			1290 => std_logic_vector(to_unsigned(228, 8)),
			1291 => std_logic_vector(to_unsigned(184, 8)),
			1292 => std_logic_vector(to_unsigned(157, 8)),
			1293 => std_logic_vector(to_unsigned(70, 8)),
			1294 => std_logic_vector(to_unsigned(35, 8)),
			1295 => std_logic_vector(to_unsigned(71, 8)),
			1296 => std_logic_vector(to_unsigned(25, 8)),
			1297 => std_logic_vector(to_unsigned(254, 8)),
			1298 => std_logic_vector(to_unsigned(45, 8)),
			1299 => std_logic_vector(to_unsigned(163, 8)),
			1300 => std_logic_vector(to_unsigned(70, 8)),
			1301 => std_logic_vector(to_unsigned(68, 8)),
			1302 => std_logic_vector(to_unsigned(57, 8)),
			1303 => std_logic_vector(to_unsigned(72, 8)),
			1304 => std_logic_vector(to_unsigned(15, 8)),
			1305 => std_logic_vector(to_unsigned(101, 8)),
			1306 => std_logic_vector(to_unsigned(86, 8)),
			1307 => std_logic_vector(to_unsigned(185, 8)),
			1308 => std_logic_vector(to_unsigned(116, 8)),
			1309 => std_logic_vector(to_unsigned(216, 8)),
			1310 => std_logic_vector(to_unsigned(209, 8)),
			1311 => std_logic_vector(to_unsigned(23, 8)),
			1312 => std_logic_vector(to_unsigned(239, 8)),
			1313 => std_logic_vector(to_unsigned(123, 8)),
			1314 => std_logic_vector(to_unsigned(216, 8)),
			1315 => std_logic_vector(to_unsigned(1, 8)),
			1316 => std_logic_vector(to_unsigned(138, 8)),
			1317 => std_logic_vector(to_unsigned(205, 8)),
			1318 => std_logic_vector(to_unsigned(167, 8)),
			1319 => std_logic_vector(to_unsigned(252, 8)),
			1320 => std_logic_vector(to_unsigned(42, 8)),
			1321 => std_logic_vector(to_unsigned(191, 8)),
			1322 => std_logic_vector(to_unsigned(3, 8)),
			1323 => std_logic_vector(to_unsigned(222, 8)),
			1324 => std_logic_vector(to_unsigned(223, 8)),
			1325 => std_logic_vector(to_unsigned(127, 8)),
			1326 => std_logic_vector(to_unsigned(0, 8)),
			1327 => std_logic_vector(to_unsigned(80, 8)),
			1328 => std_logic_vector(to_unsigned(169, 8)),
			1329 => std_logic_vector(to_unsigned(109, 8)),
			1330 => std_logic_vector(to_unsigned(187, 8)),
			1331 => std_logic_vector(to_unsigned(105, 8)),
			1332 => std_logic_vector(to_unsigned(180, 8)),
			1333 => std_logic_vector(to_unsigned(209, 8)),
			1334 => std_logic_vector(to_unsigned(187, 8)),
			1335 => std_logic_vector(to_unsigned(247, 8)),
			1336 => std_logic_vector(to_unsigned(174, 8)),
			1337 => std_logic_vector(to_unsigned(240, 8)),
			1338 => std_logic_vector(to_unsigned(156, 8)),
			1339 => std_logic_vector(to_unsigned(44, 8)),
			1340 => std_logic_vector(to_unsigned(251, 8)),
			1341 => std_logic_vector(to_unsigned(14, 8)),
			1342 => std_logic_vector(to_unsigned(224, 8)),
			1343 => std_logic_vector(to_unsigned(77, 8)),
			1344 => std_logic_vector(to_unsigned(26, 8)),
			1345 => std_logic_vector(to_unsigned(35, 8)),
			1346 => std_logic_vector(to_unsigned(18, 8)),
			1347 => std_logic_vector(to_unsigned(192, 8)),
			1348 => std_logic_vector(to_unsigned(178, 8)),
			1349 => std_logic_vector(to_unsigned(144, 8)),
			1350 => std_logic_vector(to_unsigned(43, 8)),
			1351 => std_logic_vector(to_unsigned(110, 8)),
			1352 => std_logic_vector(to_unsigned(125, 8)),
			1353 => std_logic_vector(to_unsigned(248, 8)),
			1354 => std_logic_vector(to_unsigned(33, 8)),
			1355 => std_logic_vector(to_unsigned(49, 8)),
			1356 => std_logic_vector(to_unsigned(114, 8)),
			1357 => std_logic_vector(to_unsigned(162, 8)),
			1358 => std_logic_vector(to_unsigned(56, 8)),
			1359 => std_logic_vector(to_unsigned(238, 8)),
			1360 => std_logic_vector(to_unsigned(148, 8)),
			1361 => std_logic_vector(to_unsigned(237, 8)),
			1362 => std_logic_vector(to_unsigned(157, 8)),
			1363 => std_logic_vector(to_unsigned(52, 8)),
			1364 => std_logic_vector(to_unsigned(123, 8)),
			1365 => std_logic_vector(to_unsigned(104, 8)),
			1366 => std_logic_vector(to_unsigned(141, 8)),
			1367 => std_logic_vector(to_unsigned(163, 8)),
			1368 => std_logic_vector(to_unsigned(27, 8)),
			1369 => std_logic_vector(to_unsigned(108, 8)),
			1370 => std_logic_vector(to_unsigned(174, 8)),
			1371 => std_logic_vector(to_unsigned(191, 8)),
			1372 => std_logic_vector(to_unsigned(242, 8)),
			1373 => std_logic_vector(to_unsigned(178, 8)),
			1374 => std_logic_vector(to_unsigned(14, 8)),
			1375 => std_logic_vector(to_unsigned(202, 8)),
			1376 => std_logic_vector(to_unsigned(72, 8)),
			1377 => std_logic_vector(to_unsigned(48, 8)),
			1378 => std_logic_vector(to_unsigned(83, 8)),
			1379 => std_logic_vector(to_unsigned(148, 8)),
			1380 => std_logic_vector(to_unsigned(225, 8)),
			1381 => std_logic_vector(to_unsigned(138, 8)),
			1382 => std_logic_vector(to_unsigned(235, 8)),
			1383 => std_logic_vector(to_unsigned(123, 8)),
			1384 => std_logic_vector(to_unsigned(2, 8)),
			1385 => std_logic_vector(to_unsigned(231, 8)),
			1386 => std_logic_vector(to_unsigned(7, 8)),
			1387 => std_logic_vector(to_unsigned(195, 8)),
			1388 => std_logic_vector(to_unsigned(28, 8)),
			1389 => std_logic_vector(to_unsigned(5, 8)),
			1390 => std_logic_vector(to_unsigned(179, 8)),
			1391 => std_logic_vector(to_unsigned(5, 8)),
			1392 => std_logic_vector(to_unsigned(132, 8)),
			1393 => std_logic_vector(to_unsigned(112, 8)),
			1394 => std_logic_vector(to_unsigned(93, 8)),
			1395 => std_logic_vector(to_unsigned(99, 8)),
			1396 => std_logic_vector(to_unsigned(168, 8)),
			1397 => std_logic_vector(to_unsigned(145, 8)),
			1398 => std_logic_vector(to_unsigned(70, 8)),
			1399 => std_logic_vector(to_unsigned(38, 8)),
			1400 => std_logic_vector(to_unsigned(193, 8)),
			1401 => std_logic_vector(to_unsigned(112, 8)),
			1402 => std_logic_vector(to_unsigned(213, 8)),
			1403 => std_logic_vector(to_unsigned(246, 8)),
			1404 => std_logic_vector(to_unsigned(36, 8)),
			1405 => std_logic_vector(to_unsigned(117, 8)),
			1406 => std_logic_vector(to_unsigned(135, 8)),
			1407 => std_logic_vector(to_unsigned(78, 8)),
			1408 => std_logic_vector(to_unsigned(210, 8)),
			1409 => std_logic_vector(to_unsigned(82, 8)),
			1410 => std_logic_vector(to_unsigned(18, 8)),
			1411 => std_logic_vector(to_unsigned(87, 8)),
			1412 => std_logic_vector(to_unsigned(68, 8)),
			1413 => std_logic_vector(to_unsigned(18, 8)),
			1414 => std_logic_vector(to_unsigned(50, 8)),
			1415 => std_logic_vector(to_unsigned(138, 8)),
			1416 => std_logic_vector(to_unsigned(6, 8)),
			1417 => std_logic_vector(to_unsigned(190, 8)),
			1418 => std_logic_vector(to_unsigned(200, 8)),
			1419 => std_logic_vector(to_unsigned(248, 8)),
			1420 => std_logic_vector(to_unsigned(71, 8)),
			1421 => std_logic_vector(to_unsigned(143, 8)),
			1422 => std_logic_vector(to_unsigned(127, 8)),
			1423 => std_logic_vector(to_unsigned(94, 8)),
			1424 => std_logic_vector(to_unsigned(68, 8)),
			1425 => std_logic_vector(to_unsigned(29, 8)),
			1426 => std_logic_vector(to_unsigned(155, 8)),
			1427 => std_logic_vector(to_unsigned(137, 8)),
			1428 => std_logic_vector(to_unsigned(49, 8)),
			1429 => std_logic_vector(to_unsigned(174, 8)),
			1430 => std_logic_vector(to_unsigned(104, 8)),
			1431 => std_logic_vector(to_unsigned(35, 8)),
			1432 => std_logic_vector(to_unsigned(57, 8)),
			1433 => std_logic_vector(to_unsigned(57, 8)),
			1434 => std_logic_vector(to_unsigned(74, 8)),
			1435 => std_logic_vector(to_unsigned(176, 8)),
			1436 => std_logic_vector(to_unsigned(96, 8)),
			1437 => std_logic_vector(to_unsigned(145, 8)),
			1438 => std_logic_vector(to_unsigned(109, 8)),
			1439 => std_logic_vector(to_unsigned(193, 8)),
			1440 => std_logic_vector(to_unsigned(167, 8)),
			1441 => std_logic_vector(to_unsigned(147, 8)),
			1442 => std_logic_vector(to_unsigned(78, 8)),
			1443 => std_logic_vector(to_unsigned(239, 8)),
			1444 => std_logic_vector(to_unsigned(85, 8)),
			1445 => std_logic_vector(to_unsigned(35, 8)),
			1446 => std_logic_vector(to_unsigned(255, 8)),
			1447 => std_logic_vector(to_unsigned(241, 8)),
			1448 => std_logic_vector(to_unsigned(195, 8)),
			1449 => std_logic_vector(to_unsigned(194, 8)),
			1450 => std_logic_vector(to_unsigned(209, 8)),
			1451 => std_logic_vector(to_unsigned(74, 8)),
			1452 => std_logic_vector(to_unsigned(79, 8)),
			1453 => std_logic_vector(to_unsigned(0, 8)),
			1454 => std_logic_vector(to_unsigned(210, 8)),
			1455 => std_logic_vector(to_unsigned(27, 8)),
			1456 => std_logic_vector(to_unsigned(58, 8)),
			1457 => std_logic_vector(to_unsigned(234, 8)),
			1458 => std_logic_vector(to_unsigned(220, 8)),
			1459 => std_logic_vector(to_unsigned(204, 8)),
			1460 => std_logic_vector(to_unsigned(180, 8)),
			1461 => std_logic_vector(to_unsigned(195, 8)),
			1462 => std_logic_vector(to_unsigned(94, 8)),
			1463 => std_logic_vector(to_unsigned(0, 8)),
			1464 => std_logic_vector(to_unsigned(175, 8)),
			1465 => std_logic_vector(to_unsigned(67, 8)),
			1466 => std_logic_vector(to_unsigned(246, 8)),
			1467 => std_logic_vector(to_unsigned(227, 8)),
			1468 => std_logic_vector(to_unsigned(18, 8)),
			1469 => std_logic_vector(to_unsigned(25, 8)),
			1470 => std_logic_vector(to_unsigned(155, 8)),
			1471 => std_logic_vector(to_unsigned(62, 8)),
			1472 => std_logic_vector(to_unsigned(121, 8)),
			1473 => std_logic_vector(to_unsigned(155, 8)),
			1474 => std_logic_vector(to_unsigned(23, 8)),
			1475 => std_logic_vector(to_unsigned(181, 8)),
			1476 => std_logic_vector(to_unsigned(238, 8)),
			1477 => std_logic_vector(to_unsigned(118, 8)),
			1478 => std_logic_vector(to_unsigned(5, 8)),
			1479 => std_logic_vector(to_unsigned(123, 8)),
			1480 => std_logic_vector(to_unsigned(61, 8)),
			1481 => std_logic_vector(to_unsigned(5, 8)),
			1482 => std_logic_vector(to_unsigned(86, 8)),
			1483 => std_logic_vector(to_unsigned(231, 8)),
			1484 => std_logic_vector(to_unsigned(211, 8)),
			1485 => std_logic_vector(to_unsigned(62, 8)),
			1486 => std_logic_vector(to_unsigned(80, 8)),
			1487 => std_logic_vector(to_unsigned(242, 8)),
			1488 => std_logic_vector(to_unsigned(229, 8)),
			1489 => std_logic_vector(to_unsigned(230, 8)),
			1490 => std_logic_vector(to_unsigned(160, 8)),
			1491 => std_logic_vector(to_unsigned(0, 8)),
			1492 => std_logic_vector(to_unsigned(111, 8)),
			1493 => std_logic_vector(to_unsigned(28, 8)),
			1494 => std_logic_vector(to_unsigned(173, 8)),
			1495 => std_logic_vector(to_unsigned(73, 8)),
			1496 => std_logic_vector(to_unsigned(95, 8)),
			1497 => std_logic_vector(to_unsigned(27, 8)),
			1498 => std_logic_vector(to_unsigned(215, 8)),
			1499 => std_logic_vector(to_unsigned(84, 8)),
			1500 => std_logic_vector(to_unsigned(37, 8)),
			1501 => std_logic_vector(to_unsigned(27, 8)),
			1502 => std_logic_vector(to_unsigned(94, 8)),
			1503 => std_logic_vector(to_unsigned(25, 8)),
			1504 => std_logic_vector(to_unsigned(93, 8)),
			1505 => std_logic_vector(to_unsigned(170, 8)),
			1506 => std_logic_vector(to_unsigned(163, 8)),
			1507 => std_logic_vector(to_unsigned(240, 8)),
			1508 => std_logic_vector(to_unsigned(122, 8)),
			1509 => std_logic_vector(to_unsigned(115, 8)),
			1510 => std_logic_vector(to_unsigned(107, 8)),
			1511 => std_logic_vector(to_unsigned(224, 8)),
			1512 => std_logic_vector(to_unsigned(200, 8)),
			1513 => std_logic_vector(to_unsigned(210, 8)),
			1514 => std_logic_vector(to_unsigned(57, 8)),
			1515 => std_logic_vector(to_unsigned(167, 8)),
			1516 => std_logic_vector(to_unsigned(56, 8)),
			1517 => std_logic_vector(to_unsigned(41, 8)),
			1518 => std_logic_vector(to_unsigned(225, 8)),
			1519 => std_logic_vector(to_unsigned(207, 8)),
			1520 => std_logic_vector(to_unsigned(234, 8)),
			1521 => std_logic_vector(to_unsigned(161, 8)),
			1522 => std_logic_vector(to_unsigned(7, 8)),
			1523 => std_logic_vector(to_unsigned(37, 8)),
			1524 => std_logic_vector(to_unsigned(140, 8)),
			1525 => std_logic_vector(to_unsigned(174, 8)),
			1526 => std_logic_vector(to_unsigned(102, 8)),
			1527 => std_logic_vector(to_unsigned(194, 8)),
			1528 => std_logic_vector(to_unsigned(24, 8)),
			1529 => std_logic_vector(to_unsigned(89, 8)),
			1530 => std_logic_vector(to_unsigned(170, 8)),
			1531 => std_logic_vector(to_unsigned(218, 8)),
			1532 => std_logic_vector(to_unsigned(73, 8)),
			1533 => std_logic_vector(to_unsigned(33, 8)),
			1534 => std_logic_vector(to_unsigned(1, 8)),
			1535 => std_logic_vector(to_unsigned(205, 8)),
			1536 => std_logic_vector(to_unsigned(2, 8)),
			1537 => std_logic_vector(to_unsigned(231, 8)),
			1538 => std_logic_vector(to_unsigned(147, 8)),
			1539 => std_logic_vector(to_unsigned(226, 8)),
			1540 => std_logic_vector(to_unsigned(142, 8)),
			1541 => std_logic_vector(to_unsigned(226, 8)),
			1542 => std_logic_vector(to_unsigned(12, 8)),
			1543 => std_logic_vector(to_unsigned(26, 8)),
			1544 => std_logic_vector(to_unsigned(116, 8)),
			1545 => std_logic_vector(to_unsigned(133, 8)),
			1546 => std_logic_vector(to_unsigned(64, 8)),
			1547 => std_logic_vector(to_unsigned(121, 8)),
			1548 => std_logic_vector(to_unsigned(44, 8)),
			1549 => std_logic_vector(to_unsigned(113, 8)),
			1550 => std_logic_vector(to_unsigned(127, 8)),
			1551 => std_logic_vector(to_unsigned(5, 8)),
			1552 => std_logic_vector(to_unsigned(70, 8)),
			1553 => std_logic_vector(to_unsigned(59, 8)),
			1554 => std_logic_vector(to_unsigned(233, 8)),
			1555 => std_logic_vector(to_unsigned(109, 8)),
			1556 => std_logic_vector(to_unsigned(68, 8)),
			1557 => std_logic_vector(to_unsigned(118, 8)),
			1558 => std_logic_vector(to_unsigned(173, 8)),
			1559 => std_logic_vector(to_unsigned(101, 8)),
			1560 => std_logic_vector(to_unsigned(26, 8)),
			1561 => std_logic_vector(to_unsigned(149, 8)),
			1562 => std_logic_vector(to_unsigned(255, 8)),
			1563 => std_logic_vector(to_unsigned(0, 8)),
			1564 => std_logic_vector(to_unsigned(167, 8)),
			1565 => std_logic_vector(to_unsigned(144, 8)),
			1566 => std_logic_vector(to_unsigned(44, 8)),
			1567 => std_logic_vector(to_unsigned(95, 8)),
			1568 => std_logic_vector(to_unsigned(133, 8)),
			1569 => std_logic_vector(to_unsigned(106, 8)),
			1570 => std_logic_vector(to_unsigned(209, 8)),
			1571 => std_logic_vector(to_unsigned(130, 8)),
			1572 => std_logic_vector(to_unsigned(235, 8)),
			1573 => std_logic_vector(to_unsigned(91, 8)),
			1574 => std_logic_vector(to_unsigned(86, 8)),
			1575 => std_logic_vector(to_unsigned(20, 8)),
			1576 => std_logic_vector(to_unsigned(217, 8)),
			1577 => std_logic_vector(to_unsigned(10, 8)),
			1578 => std_logic_vector(to_unsigned(59, 8)),
			1579 => std_logic_vector(to_unsigned(132, 8)),
			1580 => std_logic_vector(to_unsigned(247, 8)),
			1581 => std_logic_vector(to_unsigned(150, 8)),
			1582 => std_logic_vector(to_unsigned(204, 8)),
			1583 => std_logic_vector(to_unsigned(101, 8)),
			1584 => std_logic_vector(to_unsigned(158, 8)),
			1585 => std_logic_vector(to_unsigned(149, 8)),
			1586 => std_logic_vector(to_unsigned(211, 8)),
			1587 => std_logic_vector(to_unsigned(167, 8)),
			1588 => std_logic_vector(to_unsigned(140, 8)),
			1589 => std_logic_vector(to_unsigned(182, 8)),
			1590 => std_logic_vector(to_unsigned(165, 8)),
			1591 => std_logic_vector(to_unsigned(124, 8)),
			1592 => std_logic_vector(to_unsigned(71, 8)),
			1593 => std_logic_vector(to_unsigned(175, 8)),
			1594 => std_logic_vector(to_unsigned(137, 8)),
			1595 => std_logic_vector(to_unsigned(130, 8)),
			1596 => std_logic_vector(to_unsigned(81, 8)),
			1597 => std_logic_vector(to_unsigned(254, 8)),
			1598 => std_logic_vector(to_unsigned(65, 8)),
			1599 => std_logic_vector(to_unsigned(119, 8)),
			1600 => std_logic_vector(to_unsigned(231, 8)),
			1601 => std_logic_vector(to_unsigned(40, 8)),
			1602 => std_logic_vector(to_unsigned(208, 8)),
			1603 => std_logic_vector(to_unsigned(206, 8)),
			1604 => std_logic_vector(to_unsigned(197, 8)),
			1605 => std_logic_vector(to_unsigned(182, 8)),
			1606 => std_logic_vector(to_unsigned(130, 8)),
			1607 => std_logic_vector(to_unsigned(11, 8)),
			1608 => std_logic_vector(to_unsigned(20, 8)),
			1609 => std_logic_vector(to_unsigned(191, 8)),
			1610 => std_logic_vector(to_unsigned(9, 8)),
			1611 => std_logic_vector(to_unsigned(47, 8)),
			1612 => std_logic_vector(to_unsigned(95, 8)),
			1613 => std_logic_vector(to_unsigned(184, 8)),
			1614 => std_logic_vector(to_unsigned(142, 8)),
			1615 => std_logic_vector(to_unsigned(170, 8)),
			1616 => std_logic_vector(to_unsigned(239, 8)),
			1617 => std_logic_vector(to_unsigned(200, 8)),
			1618 => std_logic_vector(to_unsigned(60, 8)),
			1619 => std_logic_vector(to_unsigned(217, 8)),
			1620 => std_logic_vector(to_unsigned(178, 8)),
			1621 => std_logic_vector(to_unsigned(240, 8)),
			1622 => std_logic_vector(to_unsigned(10, 8)),
			1623 => std_logic_vector(to_unsigned(178, 8)),
			1624 => std_logic_vector(to_unsigned(35, 8)),
			1625 => std_logic_vector(to_unsigned(118, 8)),
			1626 => std_logic_vector(to_unsigned(28, 8)),
			1627 => std_logic_vector(to_unsigned(52, 8)),
			1628 => std_logic_vector(to_unsigned(50, 8)),
			1629 => std_logic_vector(to_unsigned(7, 8)),
			1630 => std_logic_vector(to_unsigned(153, 8)),
			1631 => std_logic_vector(to_unsigned(234, 8)),
			1632 => std_logic_vector(to_unsigned(59, 8)),
			1633 => std_logic_vector(to_unsigned(15, 8)),
			1634 => std_logic_vector(to_unsigned(226, 8)),
			1635 => std_logic_vector(to_unsigned(118, 8)),
			1636 => std_logic_vector(to_unsigned(109, 8)),
			1637 => std_logic_vector(to_unsigned(231, 8)),
			1638 => std_logic_vector(to_unsigned(187, 8)),
			1639 => std_logic_vector(to_unsigned(191, 8)),
			1640 => std_logic_vector(to_unsigned(217, 8)),
			1641 => std_logic_vector(to_unsigned(241, 8)),
			1642 => std_logic_vector(to_unsigned(156, 8)),
			1643 => std_logic_vector(to_unsigned(140, 8)),
			1644 => std_logic_vector(to_unsigned(55, 8)),
			1645 => std_logic_vector(to_unsigned(46, 8)),
			1646 => std_logic_vector(to_unsigned(196, 8)),
			1647 => std_logic_vector(to_unsigned(196, 8)),
			1648 => std_logic_vector(to_unsigned(172, 8)),
			1649 => std_logic_vector(to_unsigned(232, 8)),
			1650 => std_logic_vector(to_unsigned(255, 8)),
			1651 => std_logic_vector(to_unsigned(92, 8)),
			1652 => std_logic_vector(to_unsigned(206, 8)),
			1653 => std_logic_vector(to_unsigned(199, 8)),
			1654 => std_logic_vector(to_unsigned(211, 8)),
			1655 => std_logic_vector(to_unsigned(39, 8)),
			1656 => std_logic_vector(to_unsigned(46, 8)),
			1657 => std_logic_vector(to_unsigned(105, 8)),
			1658 => std_logic_vector(to_unsigned(145, 8)),
			1659 => std_logic_vector(to_unsigned(121, 8)),
			1660 => std_logic_vector(to_unsigned(154, 8)),
			1661 => std_logic_vector(to_unsigned(200, 8)),
			1662 => std_logic_vector(to_unsigned(130, 8)),
			1663 => std_logic_vector(to_unsigned(211, 8)),
			1664 => std_logic_vector(to_unsigned(62, 8)),
			1665 => std_logic_vector(to_unsigned(31, 8)),
			1666 => std_logic_vector(to_unsigned(35, 8)),
			1667 => std_logic_vector(to_unsigned(96, 8)),
			1668 => std_logic_vector(to_unsigned(227, 8)),
			1669 => std_logic_vector(to_unsigned(125, 8)),
			1670 => std_logic_vector(to_unsigned(195, 8)),
			1671 => std_logic_vector(to_unsigned(161, 8)),
			1672 => std_logic_vector(to_unsigned(19, 8)),
			1673 => std_logic_vector(to_unsigned(57, 8)),
			1674 => std_logic_vector(to_unsigned(131, 8)),
			1675 => std_logic_vector(to_unsigned(154, 8)),
			1676 => std_logic_vector(to_unsigned(24, 8)),
			1677 => std_logic_vector(to_unsigned(158, 8)),
			1678 => std_logic_vector(to_unsigned(78, 8)),
			1679 => std_logic_vector(to_unsigned(239, 8)),
			1680 => std_logic_vector(to_unsigned(82, 8)),
			1681 => std_logic_vector(to_unsigned(149, 8)),
			1682 => std_logic_vector(to_unsigned(73, 8)),
			1683 => std_logic_vector(to_unsigned(50, 8)),
			1684 => std_logic_vector(to_unsigned(39, 8)),
			1685 => std_logic_vector(to_unsigned(118, 8)),
			1686 => std_logic_vector(to_unsigned(19, 8)),
			1687 => std_logic_vector(to_unsigned(227, 8)),
			1688 => std_logic_vector(to_unsigned(16, 8)),
			1689 => std_logic_vector(to_unsigned(101, 8)),
			1690 => std_logic_vector(to_unsigned(20, 8)),
			1691 => std_logic_vector(to_unsigned(103, 8)),
			1692 => std_logic_vector(to_unsigned(85, 8)),
			1693 => std_logic_vector(to_unsigned(145, 8)),
			1694 => std_logic_vector(to_unsigned(242, 8)),
			1695 => std_logic_vector(to_unsigned(162, 8)),
			1696 => std_logic_vector(to_unsigned(214, 8)),
			1697 => std_logic_vector(to_unsigned(74, 8)),
			1698 => std_logic_vector(to_unsigned(49, 8)),
			1699 => std_logic_vector(to_unsigned(89, 8)),
			1700 => std_logic_vector(to_unsigned(222, 8)),
			1701 => std_logic_vector(to_unsigned(42, 8)),
			1702 => std_logic_vector(to_unsigned(35, 8)),
			1703 => std_logic_vector(to_unsigned(141, 8)),
			1704 => std_logic_vector(to_unsigned(123, 8)),
			1705 => std_logic_vector(to_unsigned(101, 8)),
			1706 => std_logic_vector(to_unsigned(213, 8)),
			1707 => std_logic_vector(to_unsigned(171, 8)),
			1708 => std_logic_vector(to_unsigned(19, 8)),
			1709 => std_logic_vector(to_unsigned(230, 8)),
			1710 => std_logic_vector(to_unsigned(211, 8)),
			1711 => std_logic_vector(to_unsigned(98, 8)),
			1712 => std_logic_vector(to_unsigned(110, 8)),
			1713 => std_logic_vector(to_unsigned(245, 8)),
			1714 => std_logic_vector(to_unsigned(247, 8)),
			1715 => std_logic_vector(to_unsigned(244, 8)),
			1716 => std_logic_vector(to_unsigned(197, 8)),
			1717 => std_logic_vector(to_unsigned(74, 8)),
			1718 => std_logic_vector(to_unsigned(127, 8)),
			1719 => std_logic_vector(to_unsigned(175, 8)),
			1720 => std_logic_vector(to_unsigned(20, 8)),
			1721 => std_logic_vector(to_unsigned(229, 8)),
			1722 => std_logic_vector(to_unsigned(210, 8)),
			1723 => std_logic_vector(to_unsigned(167, 8)),
			1724 => std_logic_vector(to_unsigned(248, 8)),
			1725 => std_logic_vector(to_unsigned(104, 8)),
			1726 => std_logic_vector(to_unsigned(7, 8)),
			1727 => std_logic_vector(to_unsigned(53, 8)),
			1728 => std_logic_vector(to_unsigned(149, 8)),
			1729 => std_logic_vector(to_unsigned(222, 8)),
			1730 => std_logic_vector(to_unsigned(251, 8)),
			1731 => std_logic_vector(to_unsigned(226, 8)),
			1732 => std_logic_vector(to_unsigned(235, 8)),
			1733 => std_logic_vector(to_unsigned(202, 8)),
			1734 => std_logic_vector(to_unsigned(229, 8)),
			1735 => std_logic_vector(to_unsigned(95, 8)),
			1736 => std_logic_vector(to_unsigned(50, 8)),
			1737 => std_logic_vector(to_unsigned(184, 8)),
			1738 => std_logic_vector(to_unsigned(171, 8)),
			1739 => std_logic_vector(to_unsigned(152, 8)),
			1740 => std_logic_vector(to_unsigned(141, 8)),
			1741 => std_logic_vector(to_unsigned(97, 8)),
			1742 => std_logic_vector(to_unsigned(139, 8)),
			1743 => std_logic_vector(to_unsigned(122, 8)),
			1744 => std_logic_vector(to_unsigned(194, 8)),
			1745 => std_logic_vector(to_unsigned(140, 8)),
			1746 => std_logic_vector(to_unsigned(157, 8)),
			1747 => std_logic_vector(to_unsigned(164, 8)),
			1748 => std_logic_vector(to_unsigned(164, 8)),
			1749 => std_logic_vector(to_unsigned(14, 8)),
			1750 => std_logic_vector(to_unsigned(194, 8)),
			1751 => std_logic_vector(to_unsigned(148, 8)),
			1752 => std_logic_vector(to_unsigned(101, 8)),
			1753 => std_logic_vector(to_unsigned(165, 8)),
			1754 => std_logic_vector(to_unsigned(206, 8)),
			1755 => std_logic_vector(to_unsigned(254, 8)),
			1756 => std_logic_vector(to_unsigned(111, 8)),
			1757 => std_logic_vector(to_unsigned(17, 8)),
			1758 => std_logic_vector(to_unsigned(135, 8)),
			1759 => std_logic_vector(to_unsigned(161, 8)),
			1760 => std_logic_vector(to_unsigned(243, 8)),
			1761 => std_logic_vector(to_unsigned(30, 8)),
			1762 => std_logic_vector(to_unsigned(82, 8)),
			1763 => std_logic_vector(to_unsigned(113, 8)),
			1764 => std_logic_vector(to_unsigned(21, 8)),
			1765 => std_logic_vector(to_unsigned(122, 8)),
			1766 => std_logic_vector(to_unsigned(14, 8)),
			1767 => std_logic_vector(to_unsigned(164, 8)),
			1768 => std_logic_vector(to_unsigned(45, 8)),
			1769 => std_logic_vector(to_unsigned(39, 8)),
			1770 => std_logic_vector(to_unsigned(149, 8)),
			1771 => std_logic_vector(to_unsigned(89, 8)),
			1772 => std_logic_vector(to_unsigned(65, 8)),
			1773 => std_logic_vector(to_unsigned(195, 8)),
			1774 => std_logic_vector(to_unsigned(201, 8)),
			1775 => std_logic_vector(to_unsigned(88, 8)),
			1776 => std_logic_vector(to_unsigned(141, 8)),
			1777 => std_logic_vector(to_unsigned(55, 8)),
			1778 => std_logic_vector(to_unsigned(190, 8)),
			1779 => std_logic_vector(to_unsigned(203, 8)),
			1780 => std_logic_vector(to_unsigned(252, 8)),
			1781 => std_logic_vector(to_unsigned(36, 8)),
			1782 => std_logic_vector(to_unsigned(14, 8)),
			1783 => std_logic_vector(to_unsigned(171, 8)),
			1784 => std_logic_vector(to_unsigned(148, 8)),
			1785 => std_logic_vector(to_unsigned(106, 8)),
			1786 => std_logic_vector(to_unsigned(193, 8)),
			1787 => std_logic_vector(to_unsigned(222, 8)),
			1788 => std_logic_vector(to_unsigned(180, 8)),
			1789 => std_logic_vector(to_unsigned(113, 8)),
			1790 => std_logic_vector(to_unsigned(253, 8)),
			1791 => std_logic_vector(to_unsigned(54, 8)),
			1792 => std_logic_vector(to_unsigned(4, 8)),
			1793 => std_logic_vector(to_unsigned(168, 8)),
			1794 => std_logic_vector(to_unsigned(13, 8)),
			1795 => std_logic_vector(to_unsigned(58, 8)),
			1796 => std_logic_vector(to_unsigned(61, 8)),
			1797 => std_logic_vector(to_unsigned(75, 8)),
			1798 => std_logic_vector(to_unsigned(30, 8)),
			1799 => std_logic_vector(to_unsigned(120, 8)),
			1800 => std_logic_vector(to_unsigned(11, 8)),
			1801 => std_logic_vector(to_unsigned(239, 8)),
			1802 => std_logic_vector(to_unsigned(49, 8)),
			1803 => std_logic_vector(to_unsigned(250, 8)),
			1804 => std_logic_vector(to_unsigned(254, 8)),
			1805 => std_logic_vector(to_unsigned(214, 8)),
			1806 => std_logic_vector(to_unsigned(3, 8)),
			1807 => std_logic_vector(to_unsigned(150, 8)),
			1808 => std_logic_vector(to_unsigned(72, 8)),
			1809 => std_logic_vector(to_unsigned(151, 8)),
			1810 => std_logic_vector(to_unsigned(115, 8)),
			1811 => std_logic_vector(to_unsigned(48, 8)),
			1812 => std_logic_vector(to_unsigned(219, 8)),
			1813 => std_logic_vector(to_unsigned(171, 8)),
			1814 => std_logic_vector(to_unsigned(119, 8)),
			1815 => std_logic_vector(to_unsigned(152, 8)),
			1816 => std_logic_vector(to_unsigned(177, 8)),
			1817 => std_logic_vector(to_unsigned(4, 8)),
			1818 => std_logic_vector(to_unsigned(73, 8)),
			1819 => std_logic_vector(to_unsigned(135, 8)),
			1820 => std_logic_vector(to_unsigned(237, 8)),
			1821 => std_logic_vector(to_unsigned(138, 8)),
			1822 => std_logic_vector(to_unsigned(204, 8)),
			1823 => std_logic_vector(to_unsigned(173, 8)),
			1824 => std_logic_vector(to_unsigned(13, 8)),
			1825 => std_logic_vector(to_unsigned(67, 8)),
			1826 => std_logic_vector(to_unsigned(57, 8)),
			1827 => std_logic_vector(to_unsigned(92, 8)),
			1828 => std_logic_vector(to_unsigned(229, 8)),
			1829 => std_logic_vector(to_unsigned(191, 8)),
			1830 => std_logic_vector(to_unsigned(125, 8)),
			1831 => std_logic_vector(to_unsigned(156, 8)),
			1832 => std_logic_vector(to_unsigned(16, 8)),
			1833 => std_logic_vector(to_unsigned(206, 8)),
			1834 => std_logic_vector(to_unsigned(130, 8)),
			1835 => std_logic_vector(to_unsigned(20, 8)),
			1836 => std_logic_vector(to_unsigned(179, 8)),
			1837 => std_logic_vector(to_unsigned(241, 8)),
			1838 => std_logic_vector(to_unsigned(11, 8)),
			1839 => std_logic_vector(to_unsigned(39, 8)),
			1840 => std_logic_vector(to_unsigned(218, 8)),
			1841 => std_logic_vector(to_unsigned(217, 8)),
			1842 => std_logic_vector(to_unsigned(131, 8)),
			1843 => std_logic_vector(to_unsigned(229, 8)),
			1844 => std_logic_vector(to_unsigned(79, 8)),
			1845 => std_logic_vector(to_unsigned(183, 8)),
			1846 => std_logic_vector(to_unsigned(195, 8)),
			1847 => std_logic_vector(to_unsigned(113, 8)),
			1848 => std_logic_vector(to_unsigned(201, 8)),
			1849 => std_logic_vector(to_unsigned(25, 8)),
			1850 => std_logic_vector(to_unsigned(189, 8)),
			1851 => std_logic_vector(to_unsigned(157, 8)),
			1852 => std_logic_vector(to_unsigned(63, 8)),
			1853 => std_logic_vector(to_unsigned(163, 8)),
			1854 => std_logic_vector(to_unsigned(173, 8)),
			1855 => std_logic_vector(to_unsigned(208, 8)),
			1856 => std_logic_vector(to_unsigned(82, 8)),
			1857 => std_logic_vector(to_unsigned(231, 8)),
			1858 => std_logic_vector(to_unsigned(240, 8)),
			1859 => std_logic_vector(to_unsigned(117, 8)),
			1860 => std_logic_vector(to_unsigned(114, 8)),
			1861 => std_logic_vector(to_unsigned(145, 8)),
			1862 => std_logic_vector(to_unsigned(117, 8)),
			1863 => std_logic_vector(to_unsigned(146, 8)),
			1864 => std_logic_vector(to_unsigned(214, 8)),
			1865 => std_logic_vector(to_unsigned(28, 8)),
			1866 => std_logic_vector(to_unsigned(177, 8)),
			1867 => std_logic_vector(to_unsigned(55, 8)),
			1868 => std_logic_vector(to_unsigned(1, 8)),
			1869 => std_logic_vector(to_unsigned(120, 8)),
			1870 => std_logic_vector(to_unsigned(178, 8)),
			1871 => std_logic_vector(to_unsigned(58, 8)),
			1872 => std_logic_vector(to_unsigned(134, 8)),
			1873 => std_logic_vector(to_unsigned(53, 8)),
			1874 => std_logic_vector(to_unsigned(233, 8)),
			1875 => std_logic_vector(to_unsigned(129, 8)),
			1876 => std_logic_vector(to_unsigned(159, 8)),
			1877 => std_logic_vector(to_unsigned(201, 8)),
			1878 => std_logic_vector(to_unsigned(152, 8)),
			1879 => std_logic_vector(to_unsigned(234, 8)),
			1880 => std_logic_vector(to_unsigned(188, 8)),
			1881 => std_logic_vector(to_unsigned(172, 8)),
			1882 => std_logic_vector(to_unsigned(28, 8)),
			1883 => std_logic_vector(to_unsigned(31, 8)),
			1884 => std_logic_vector(to_unsigned(152, 8)),
			1885 => std_logic_vector(to_unsigned(86, 8)),
			1886 => std_logic_vector(to_unsigned(243, 8)),
			1887 => std_logic_vector(to_unsigned(83, 8)),
			1888 => std_logic_vector(to_unsigned(0, 8)),
			1889 => std_logic_vector(to_unsigned(96, 8)),
			1890 => std_logic_vector(to_unsigned(130, 8)),
			1891 => std_logic_vector(to_unsigned(35, 8)),
			1892 => std_logic_vector(to_unsigned(215, 8)),
			1893 => std_logic_vector(to_unsigned(109, 8)),
			1894 => std_logic_vector(to_unsigned(199, 8)),
			1895 => std_logic_vector(to_unsigned(113, 8)),
			1896 => std_logic_vector(to_unsigned(47, 8)),
			1897 => std_logic_vector(to_unsigned(152, 8)),
			1898 => std_logic_vector(to_unsigned(166, 8)),
			1899 => std_logic_vector(to_unsigned(175, 8)),
			1900 => std_logic_vector(to_unsigned(108, 8)),
			1901 => std_logic_vector(to_unsigned(174, 8)),
			1902 => std_logic_vector(to_unsigned(6, 8)),
			1903 => std_logic_vector(to_unsigned(44, 8)),
			1904 => std_logic_vector(to_unsigned(201, 8)),
			1905 => std_logic_vector(to_unsigned(208, 8)),
			1906 => std_logic_vector(to_unsigned(206, 8)),
			1907 => std_logic_vector(to_unsigned(196, 8)),
			1908 => std_logic_vector(to_unsigned(172, 8)),
			1909 => std_logic_vector(to_unsigned(116, 8)),
			1910 => std_logic_vector(to_unsigned(202, 8)),
			1911 => std_logic_vector(to_unsigned(221, 8)),
			1912 => std_logic_vector(to_unsigned(87, 8)),
			1913 => std_logic_vector(to_unsigned(158, 8)),
			1914 => std_logic_vector(to_unsigned(73, 8)),
			1915 => std_logic_vector(to_unsigned(15, 8)),
			1916 => std_logic_vector(to_unsigned(62, 8)),
			1917 => std_logic_vector(to_unsigned(105, 8)),
			1918 => std_logic_vector(to_unsigned(184, 8)),
			1919 => std_logic_vector(to_unsigned(1, 8)),
			1920 => std_logic_vector(to_unsigned(108, 8)),
			1921 => std_logic_vector(to_unsigned(255, 8)),
			1922 => std_logic_vector(to_unsigned(169, 8)),
			1923 => std_logic_vector(to_unsigned(245, 8)),
			1924 => std_logic_vector(to_unsigned(167, 8)),
			1925 => std_logic_vector(to_unsigned(226, 8)),
			1926 => std_logic_vector(to_unsigned(223, 8)),
			1927 => std_logic_vector(to_unsigned(53, 8)),
			1928 => std_logic_vector(to_unsigned(241, 8)),
			1929 => std_logic_vector(to_unsigned(153, 8)),
			1930 => std_logic_vector(to_unsigned(167, 8)),
			1931 => std_logic_vector(to_unsigned(44, 8)),
			1932 => std_logic_vector(to_unsigned(154, 8)),
			1933 => std_logic_vector(to_unsigned(205, 8)),
			1934 => std_logic_vector(to_unsigned(18, 8)),
			1935 => std_logic_vector(to_unsigned(79, 8)),
			1936 => std_logic_vector(to_unsigned(191, 8)),
			1937 => std_logic_vector(to_unsigned(216, 8)),
			1938 => std_logic_vector(to_unsigned(253, 8)),
			1939 => std_logic_vector(to_unsigned(128, 8)),
			1940 => std_logic_vector(to_unsigned(215, 8)),
			1941 => std_logic_vector(to_unsigned(143, 8)),
			1942 => std_logic_vector(to_unsigned(227, 8)),
			1943 => std_logic_vector(to_unsigned(245, 8)),
			1944 => std_logic_vector(to_unsigned(153, 8)),
			1945 => std_logic_vector(to_unsigned(40, 8)),
			1946 => std_logic_vector(to_unsigned(2, 8)),
			1947 => std_logic_vector(to_unsigned(34, 8)),
			1948 => std_logic_vector(to_unsigned(106, 8)),
			1949 => std_logic_vector(to_unsigned(215, 8)),
			1950 => std_logic_vector(to_unsigned(28, 8)),
			1951 => std_logic_vector(to_unsigned(166, 8)),
			1952 => std_logic_vector(to_unsigned(203, 8)),
			1953 => std_logic_vector(to_unsigned(31, 8)),
			1954 => std_logic_vector(to_unsigned(53, 8)),
			1955 => std_logic_vector(to_unsigned(22, 8)),
			1956 => std_logic_vector(to_unsigned(231, 8)),
			1957 => std_logic_vector(to_unsigned(128, 8)),
			1958 => std_logic_vector(to_unsigned(119, 8)),
			1959 => std_logic_vector(to_unsigned(171, 8)),
			1960 => std_logic_vector(to_unsigned(63, 8)),
			1961 => std_logic_vector(to_unsigned(78, 8)),
			1962 => std_logic_vector(to_unsigned(13, 8)),
			1963 => std_logic_vector(to_unsigned(222, 8)),
			1964 => std_logic_vector(to_unsigned(179, 8)),
			1965 => std_logic_vector(to_unsigned(203, 8)),
			1966 => std_logic_vector(to_unsigned(104, 8)),
			1967 => std_logic_vector(to_unsigned(165, 8)),
			1968 => std_logic_vector(to_unsigned(216, 8)),
			1969 => std_logic_vector(to_unsigned(196, 8)),
			1970 => std_logic_vector(to_unsigned(252, 8)),
			1971 => std_logic_vector(to_unsigned(151, 8)),
			1972 => std_logic_vector(to_unsigned(37, 8)),
			1973 => std_logic_vector(to_unsigned(38, 8)),
			1974 => std_logic_vector(to_unsigned(225, 8)),
			1975 => std_logic_vector(to_unsigned(103, 8)),
			1976 => std_logic_vector(to_unsigned(244, 8)),
			1977 => std_logic_vector(to_unsigned(234, 8)),
			1978 => std_logic_vector(to_unsigned(97, 8)),
			1979 => std_logic_vector(to_unsigned(154, 8)),
			1980 => std_logic_vector(to_unsigned(248, 8)),
			1981 => std_logic_vector(to_unsigned(219, 8)),
			1982 => std_logic_vector(to_unsigned(130, 8)),
			1983 => std_logic_vector(to_unsigned(11, 8)),
			1984 => std_logic_vector(to_unsigned(50, 8)),
			1985 => std_logic_vector(to_unsigned(166, 8)),
			1986 => std_logic_vector(to_unsigned(24, 8)),
			1987 => std_logic_vector(to_unsigned(12, 8)),
			1988 => std_logic_vector(to_unsigned(187, 8)),
			1989 => std_logic_vector(to_unsigned(79, 8)),
			1990 => std_logic_vector(to_unsigned(97, 8)),
			1991 => std_logic_vector(to_unsigned(27, 8)),
			1992 => std_logic_vector(to_unsigned(180, 8)),
			1993 => std_logic_vector(to_unsigned(55, 8)),
			1994 => std_logic_vector(to_unsigned(153, 8)),
			1995 => std_logic_vector(to_unsigned(130, 8)),
			1996 => std_logic_vector(to_unsigned(191, 8)),
			1997 => std_logic_vector(to_unsigned(155, 8)),
			1998 => std_logic_vector(to_unsigned(98, 8)),
			1999 => std_logic_vector(to_unsigned(155, 8)),
			2000 => std_logic_vector(to_unsigned(154, 8)),
			2001 => std_logic_vector(to_unsigned(3, 8)),
			2002 => std_logic_vector(to_unsigned(67, 8)),
			2003 => std_logic_vector(to_unsigned(155, 8)),
			2004 => std_logic_vector(to_unsigned(233, 8)),
			2005 => std_logic_vector(to_unsigned(91, 8)),
			2006 => std_logic_vector(to_unsigned(200, 8)),
			2007 => std_logic_vector(to_unsigned(132, 8)),
			2008 => std_logic_vector(to_unsigned(67, 8)),
			2009 => std_logic_vector(to_unsigned(172, 8)),
			2010 => std_logic_vector(to_unsigned(236, 8)),
			2011 => std_logic_vector(to_unsigned(68, 8)),
			2012 => std_logic_vector(to_unsigned(54, 8)),
			2013 => std_logic_vector(to_unsigned(152, 8)),
			2014 => std_logic_vector(to_unsigned(30, 8)),
			2015 => std_logic_vector(to_unsigned(147, 8)),
			2016 => std_logic_vector(to_unsigned(253, 8)),
			2017 => std_logic_vector(to_unsigned(190, 8)),
			2018 => std_logic_vector(to_unsigned(1, 8)),
			2019 => std_logic_vector(to_unsigned(212, 8)),
			2020 => std_logic_vector(to_unsigned(132, 8)),
			2021 => std_logic_vector(to_unsigned(163, 8)),
			2022 => std_logic_vector(to_unsigned(142, 8)),
			2023 => std_logic_vector(to_unsigned(131, 8)),
			2024 => std_logic_vector(to_unsigned(254, 8)),
			2025 => std_logic_vector(to_unsigned(154, 8)),
			2026 => std_logic_vector(to_unsigned(178, 8)),
			2027 => std_logic_vector(to_unsigned(149, 8)),
			2028 => std_logic_vector(to_unsigned(21, 8)),
			2029 => std_logic_vector(to_unsigned(96, 8)),
			2030 => std_logic_vector(to_unsigned(184, 8)),
			2031 => std_logic_vector(to_unsigned(114, 8)),
			2032 => std_logic_vector(to_unsigned(85, 8)),
			2033 => std_logic_vector(to_unsigned(254, 8)),
			2034 => std_logic_vector(to_unsigned(150, 8)),
			2035 => std_logic_vector(to_unsigned(157, 8)),
			2036 => std_logic_vector(to_unsigned(228, 8)),
			2037 => std_logic_vector(to_unsigned(221, 8)),
			2038 => std_logic_vector(to_unsigned(33, 8)),
			2039 => std_logic_vector(to_unsigned(70, 8)),
			2040 => std_logic_vector(to_unsigned(42, 8)),
			2041 => std_logic_vector(to_unsigned(181, 8)),
			2042 => std_logic_vector(to_unsigned(117, 8)),
			2043 => std_logic_vector(to_unsigned(193, 8)),
			2044 => std_logic_vector(to_unsigned(215, 8)),
			2045 => std_logic_vector(to_unsigned(61, 8)),
			2046 => std_logic_vector(to_unsigned(247, 8)),
			2047 => std_logic_vector(to_unsigned(126, 8)),
			2048 => std_logic_vector(to_unsigned(9, 8)),
			2049 => std_logic_vector(to_unsigned(154, 8)),
			2050 => std_logic_vector(to_unsigned(90, 8)),
			2051 => std_logic_vector(to_unsigned(234, 8)),
			2052 => std_logic_vector(to_unsigned(37, 8)),
			2053 => std_logic_vector(to_unsigned(86, 8)),
			2054 => std_logic_vector(to_unsigned(234, 8)),
			2055 => std_logic_vector(to_unsigned(237, 8)),
			2056 => std_logic_vector(to_unsigned(181, 8)),
			2057 => std_logic_vector(to_unsigned(216, 8)),
			2058 => std_logic_vector(to_unsigned(35, 8)),
			2059 => std_logic_vector(to_unsigned(222, 8)),
			2060 => std_logic_vector(to_unsigned(100, 8)),
			2061 => std_logic_vector(to_unsigned(20, 8)),
			2062 => std_logic_vector(to_unsigned(73, 8)),
			2063 => std_logic_vector(to_unsigned(12, 8)),
			2064 => std_logic_vector(to_unsigned(185, 8)),
			2065 => std_logic_vector(to_unsigned(26, 8)),
			2066 => std_logic_vector(to_unsigned(166, 8)),
			2067 => std_logic_vector(to_unsigned(55, 8)),
			2068 => std_logic_vector(to_unsigned(249, 8)),
			2069 => std_logic_vector(to_unsigned(88, 8)),
			2070 => std_logic_vector(to_unsigned(2, 8)),
			2071 => std_logic_vector(to_unsigned(207, 8)),
			2072 => std_logic_vector(to_unsigned(203, 8)),
			2073 => std_logic_vector(to_unsigned(29, 8)),
			2074 => std_logic_vector(to_unsigned(7, 8)),
			2075 => std_logic_vector(to_unsigned(236, 8)),
			2076 => std_logic_vector(to_unsigned(247, 8)),
			2077 => std_logic_vector(to_unsigned(84, 8)),
			2078 => std_logic_vector(to_unsigned(152, 8)),
			2079 => std_logic_vector(to_unsigned(175, 8)),
			2080 => std_logic_vector(to_unsigned(99, 8)),
			2081 => std_logic_vector(to_unsigned(81, 8)),
			2082 => std_logic_vector(to_unsigned(102, 8)),
			2083 => std_logic_vector(to_unsigned(17, 8)),
			2084 => std_logic_vector(to_unsigned(255, 8)),
			2085 => std_logic_vector(to_unsigned(174, 8)),
			2086 => std_logic_vector(to_unsigned(122, 8)),
			2087 => std_logic_vector(to_unsigned(19, 8)),
			2088 => std_logic_vector(to_unsigned(58, 8)),
			2089 => std_logic_vector(to_unsigned(53, 8)),
			2090 => std_logic_vector(to_unsigned(178, 8)),
			2091 => std_logic_vector(to_unsigned(222, 8)),
			2092 => std_logic_vector(to_unsigned(20, 8)),
			2093 => std_logic_vector(to_unsigned(76, 8)),
			2094 => std_logic_vector(to_unsigned(231, 8)),
			2095 => std_logic_vector(to_unsigned(235, 8)),
			2096 => std_logic_vector(to_unsigned(69, 8)),
			2097 => std_logic_vector(to_unsigned(151, 8)),
			2098 => std_logic_vector(to_unsigned(69, 8)),
			2099 => std_logic_vector(to_unsigned(5, 8)),
			2100 => std_logic_vector(to_unsigned(25, 8)),
			2101 => std_logic_vector(to_unsigned(232, 8)),
			2102 => std_logic_vector(to_unsigned(200, 8)),
			2103 => std_logic_vector(to_unsigned(230, 8)),
			2104 => std_logic_vector(to_unsigned(30, 8)),
			2105 => std_logic_vector(to_unsigned(6, 8)),
			2106 => std_logic_vector(to_unsigned(72, 8)),
			2107 => std_logic_vector(to_unsigned(120, 8)),
			2108 => std_logic_vector(to_unsigned(48, 8)),
			2109 => std_logic_vector(to_unsigned(70, 8)),
			2110 => std_logic_vector(to_unsigned(12, 8)),
			2111 => std_logic_vector(to_unsigned(177, 8)),
			2112 => std_logic_vector(to_unsigned(185, 8)),
			2113 => std_logic_vector(to_unsigned(68, 8)),
			2114 => std_logic_vector(to_unsigned(219, 8)),
			2115 => std_logic_vector(to_unsigned(7, 8)),
			2116 => std_logic_vector(to_unsigned(24, 8)),
			2117 => std_logic_vector(to_unsigned(189, 8)),
			2118 => std_logic_vector(to_unsigned(65, 8)),
			2119 => std_logic_vector(to_unsigned(205, 8)),
			2120 => std_logic_vector(to_unsigned(182, 8)),
			2121 => std_logic_vector(to_unsigned(67, 8)),
			2122 => std_logic_vector(to_unsigned(36, 8)),
			2123 => std_logic_vector(to_unsigned(132, 8)),
			2124 => std_logic_vector(to_unsigned(147, 8)),
			2125 => std_logic_vector(to_unsigned(250, 8)),
			2126 => std_logic_vector(to_unsigned(118, 8)),
			2127 => std_logic_vector(to_unsigned(120, 8)),
			2128 => std_logic_vector(to_unsigned(105, 8)),
			2129 => std_logic_vector(to_unsigned(197, 8)),
			2130 => std_logic_vector(to_unsigned(106, 8)),
			2131 => std_logic_vector(to_unsigned(30, 8)),
			2132 => std_logic_vector(to_unsigned(116, 8)),
			2133 => std_logic_vector(to_unsigned(169, 8)),
			2134 => std_logic_vector(to_unsigned(156, 8)),
			2135 => std_logic_vector(to_unsigned(9, 8)),
			2136 => std_logic_vector(to_unsigned(158, 8)),
			2137 => std_logic_vector(to_unsigned(47, 8)),
			2138 => std_logic_vector(to_unsigned(191, 8)),
			2139 => std_logic_vector(to_unsigned(76, 8)),
			2140 => std_logic_vector(to_unsigned(203, 8)),
			2141 => std_logic_vector(to_unsigned(106, 8)),
			2142 => std_logic_vector(to_unsigned(0, 8)),
			2143 => std_logic_vector(to_unsigned(9, 8)),
			2144 => std_logic_vector(to_unsigned(225, 8)),
			2145 => std_logic_vector(to_unsigned(205, 8)),
			2146 => std_logic_vector(to_unsigned(118, 8)),
			2147 => std_logic_vector(to_unsigned(181, 8)),
			2148 => std_logic_vector(to_unsigned(95, 8)),
			2149 => std_logic_vector(to_unsigned(211, 8)),
			2150 => std_logic_vector(to_unsigned(152, 8)),
			2151 => std_logic_vector(to_unsigned(246, 8)),
			2152 => std_logic_vector(to_unsigned(34, 8)),
			2153 => std_logic_vector(to_unsigned(116, 8)),
			2154 => std_logic_vector(to_unsigned(255, 8)),
			2155 => std_logic_vector(to_unsigned(189, 8)),
			2156 => std_logic_vector(to_unsigned(120, 8)),
			2157 => std_logic_vector(to_unsigned(233, 8)),
			2158 => std_logic_vector(to_unsigned(25, 8)),
			2159 => std_logic_vector(to_unsigned(46, 8)),
			2160 => std_logic_vector(to_unsigned(152, 8)),
			2161 => std_logic_vector(to_unsigned(6, 8)),
			2162 => std_logic_vector(to_unsigned(136, 8)),
			2163 => std_logic_vector(to_unsigned(231, 8)),
			2164 => std_logic_vector(to_unsigned(234, 8)),
			2165 => std_logic_vector(to_unsigned(158, 8)),
			2166 => std_logic_vector(to_unsigned(142, 8)),
			2167 => std_logic_vector(to_unsigned(173, 8)),
			2168 => std_logic_vector(to_unsigned(254, 8)),
			2169 => std_logic_vector(to_unsigned(70, 8)),
			2170 => std_logic_vector(to_unsigned(181, 8)),
			2171 => std_logic_vector(to_unsigned(64, 8)),
			2172 => std_logic_vector(to_unsigned(4, 8)),
			2173 => std_logic_vector(to_unsigned(102, 8)),
			2174 => std_logic_vector(to_unsigned(42, 8)),
			2175 => std_logic_vector(to_unsigned(117, 8)),
			2176 => std_logic_vector(to_unsigned(14, 8)),
			2177 => std_logic_vector(to_unsigned(30, 8)),
			2178 => std_logic_vector(to_unsigned(136, 8)),
			2179 => std_logic_vector(to_unsigned(175, 8)),
			2180 => std_logic_vector(to_unsigned(189, 8)),
			2181 => std_logic_vector(to_unsigned(84, 8)),
			2182 => std_logic_vector(to_unsigned(226, 8)),
			2183 => std_logic_vector(to_unsigned(21, 8)),
			2184 => std_logic_vector(to_unsigned(81, 8)),
			2185 => std_logic_vector(to_unsigned(90, 8)),
			2186 => std_logic_vector(to_unsigned(96, 8)),
			2187 => std_logic_vector(to_unsigned(34, 8)),
			2188 => std_logic_vector(to_unsigned(255, 8)),
			2189 => std_logic_vector(to_unsigned(11, 8)),
			2190 => std_logic_vector(to_unsigned(133, 8)),
			2191 => std_logic_vector(to_unsigned(58, 8)),
			2192 => std_logic_vector(to_unsigned(172, 8)),
			2193 => std_logic_vector(to_unsigned(192, 8)),
			2194 => std_logic_vector(to_unsigned(165, 8)),
			2195 => std_logic_vector(to_unsigned(216, 8)),
			2196 => std_logic_vector(to_unsigned(219, 8)),
			2197 => std_logic_vector(to_unsigned(229, 8)),
			2198 => std_logic_vector(to_unsigned(170, 8)),
			2199 => std_logic_vector(to_unsigned(11, 8)),
			2200 => std_logic_vector(to_unsigned(221, 8)),
			2201 => std_logic_vector(to_unsigned(32, 8)),
			2202 => std_logic_vector(to_unsigned(71, 8)),
			2203 => std_logic_vector(to_unsigned(239, 8)),
			2204 => std_logic_vector(to_unsigned(245, 8)),
			2205 => std_logic_vector(to_unsigned(228, 8)),
			2206 => std_logic_vector(to_unsigned(115, 8)),
			2207 => std_logic_vector(to_unsigned(14, 8)),
			2208 => std_logic_vector(to_unsigned(208, 8)),
			2209 => std_logic_vector(to_unsigned(100, 8)),
			2210 => std_logic_vector(to_unsigned(80, 8)),
			2211 => std_logic_vector(to_unsigned(76, 8)),
			2212 => std_logic_vector(to_unsigned(200, 8)),
			2213 => std_logic_vector(to_unsigned(36, 8)),
			2214 => std_logic_vector(to_unsigned(166, 8)),
			2215 => std_logic_vector(to_unsigned(61, 8)),
			2216 => std_logic_vector(to_unsigned(135, 8)),
			2217 => std_logic_vector(to_unsigned(174, 8)),
			2218 => std_logic_vector(to_unsigned(90, 8)),
			2219 => std_logic_vector(to_unsigned(159, 8)),
			2220 => std_logic_vector(to_unsigned(135, 8)),
			2221 => std_logic_vector(to_unsigned(34, 8)),
			2222 => std_logic_vector(to_unsigned(112, 8)),
			2223 => std_logic_vector(to_unsigned(252, 8)),
			2224 => std_logic_vector(to_unsigned(245, 8)),
			2225 => std_logic_vector(to_unsigned(118, 8)),
			2226 => std_logic_vector(to_unsigned(164, 8)),
			2227 => std_logic_vector(to_unsigned(148, 8)),
			2228 => std_logic_vector(to_unsigned(21, 8)),
			2229 => std_logic_vector(to_unsigned(166, 8)),
			2230 => std_logic_vector(to_unsigned(116, 8)),
			2231 => std_logic_vector(to_unsigned(248, 8)),
			2232 => std_logic_vector(to_unsigned(118, 8)),
			2233 => std_logic_vector(to_unsigned(30, 8)),
			2234 => std_logic_vector(to_unsigned(94, 8)),
			2235 => std_logic_vector(to_unsigned(243, 8)),
			2236 => std_logic_vector(to_unsigned(193, 8)),
			2237 => std_logic_vector(to_unsigned(137, 8)),
			2238 => std_logic_vector(to_unsigned(208, 8)),
			2239 => std_logic_vector(to_unsigned(140, 8)),
			2240 => std_logic_vector(to_unsigned(148, 8)),
			2241 => std_logic_vector(to_unsigned(236, 8)),
			2242 => std_logic_vector(to_unsigned(100, 8)),
			2243 => std_logic_vector(to_unsigned(232, 8)),
			2244 => std_logic_vector(to_unsigned(100, 8)),
			2245 => std_logic_vector(to_unsigned(22, 8)),
			2246 => std_logic_vector(to_unsigned(128, 8)),
			2247 => std_logic_vector(to_unsigned(221, 8)),
			2248 => std_logic_vector(to_unsigned(66, 8)),
			2249 => std_logic_vector(to_unsigned(219, 8)),
			2250 => std_logic_vector(to_unsigned(106, 8)),
			2251 => std_logic_vector(to_unsigned(111, 8)),
			2252 => std_logic_vector(to_unsigned(232, 8)),
			2253 => std_logic_vector(to_unsigned(219, 8)),
			2254 => std_logic_vector(to_unsigned(198, 8)),
			2255 => std_logic_vector(to_unsigned(83, 8)),
			2256 => std_logic_vector(to_unsigned(70, 8)),
			2257 => std_logic_vector(to_unsigned(0, 8)),
			2258 => std_logic_vector(to_unsigned(210, 8)),
			2259 => std_logic_vector(to_unsigned(139, 8)),
			2260 => std_logic_vector(to_unsigned(124, 8)),
			2261 => std_logic_vector(to_unsigned(107, 8)),
			2262 => std_logic_vector(to_unsigned(154, 8)),
			2263 => std_logic_vector(to_unsigned(177, 8)),
			2264 => std_logic_vector(to_unsigned(26, 8)),
			2265 => std_logic_vector(to_unsigned(100, 8)),
			2266 => std_logic_vector(to_unsigned(216, 8)),
			2267 => std_logic_vector(to_unsigned(10, 8)),
			2268 => std_logic_vector(to_unsigned(206, 8)),
			2269 => std_logic_vector(to_unsigned(62, 8)),
			2270 => std_logic_vector(to_unsigned(70, 8)),
			2271 => std_logic_vector(to_unsigned(15, 8)),
			2272 => std_logic_vector(to_unsigned(161, 8)),
			2273 => std_logic_vector(to_unsigned(79, 8)),
			2274 => std_logic_vector(to_unsigned(53, 8)),
			2275 => std_logic_vector(to_unsigned(244, 8)),
			2276 => std_logic_vector(to_unsigned(12, 8)),
			2277 => std_logic_vector(to_unsigned(120, 8)),
			2278 => std_logic_vector(to_unsigned(113, 8)),
			2279 => std_logic_vector(to_unsigned(222, 8)),
			2280 => std_logic_vector(to_unsigned(116, 8)),
			2281 => std_logic_vector(to_unsigned(12, 8)),
			2282 => std_logic_vector(to_unsigned(159, 8)),
			2283 => std_logic_vector(to_unsigned(11, 8)),
			2284 => std_logic_vector(to_unsigned(4, 8)),
			2285 => std_logic_vector(to_unsigned(5, 8)),
			2286 => std_logic_vector(to_unsigned(108, 8)),
			2287 => std_logic_vector(to_unsigned(209, 8)),
			2288 => std_logic_vector(to_unsigned(3, 8)),
			2289 => std_logic_vector(to_unsigned(210, 8)),
			2290 => std_logic_vector(to_unsigned(54, 8)),
			2291 => std_logic_vector(to_unsigned(169, 8)),
			2292 => std_logic_vector(to_unsigned(180, 8)),
			2293 => std_logic_vector(to_unsigned(223, 8)),
			2294 => std_logic_vector(to_unsigned(117, 8)),
			2295 => std_logic_vector(to_unsigned(93, 8)),
			2296 => std_logic_vector(to_unsigned(142, 8)),
			2297 => std_logic_vector(to_unsigned(174, 8)),
			2298 => std_logic_vector(to_unsigned(188, 8)),
			2299 => std_logic_vector(to_unsigned(56, 8)),
			2300 => std_logic_vector(to_unsigned(160, 8)),
			2301 => std_logic_vector(to_unsigned(130, 8)),
			2302 => std_logic_vector(to_unsigned(200, 8)),
			2303 => std_logic_vector(to_unsigned(141, 8)),
			2304 => std_logic_vector(to_unsigned(242, 8)),
			2305 => std_logic_vector(to_unsigned(163, 8)),
			2306 => std_logic_vector(to_unsigned(122, 8)),
			2307 => std_logic_vector(to_unsigned(23, 8)),
			2308 => std_logic_vector(to_unsigned(255, 8)),
			2309 => std_logic_vector(to_unsigned(211, 8)),
			2310 => std_logic_vector(to_unsigned(251, 8)),
			2311 => std_logic_vector(to_unsigned(92, 8)),
			2312 => std_logic_vector(to_unsigned(120, 8)),
			2313 => std_logic_vector(to_unsigned(202, 8)),
			2314 => std_logic_vector(to_unsigned(27, 8)),
			2315 => std_logic_vector(to_unsigned(96, 8)),
			2316 => std_logic_vector(to_unsigned(46, 8)),
			2317 => std_logic_vector(to_unsigned(192, 8)),
			2318 => std_logic_vector(to_unsigned(247, 8)),
			2319 => std_logic_vector(to_unsigned(5, 8)),
			2320 => std_logic_vector(to_unsigned(227, 8)),
			2321 => std_logic_vector(to_unsigned(101, 8)),
			2322 => std_logic_vector(to_unsigned(91, 8)),
			2323 => std_logic_vector(to_unsigned(229, 8)),
			2324 => std_logic_vector(to_unsigned(2, 8)),
			2325 => std_logic_vector(to_unsigned(116, 8)),
			2326 => std_logic_vector(to_unsigned(152, 8)),
			2327 => std_logic_vector(to_unsigned(23, 8)),
			2328 => std_logic_vector(to_unsigned(205, 8)),
			2329 => std_logic_vector(to_unsigned(100, 8)),
			2330 => std_logic_vector(to_unsigned(201, 8)),
			2331 => std_logic_vector(to_unsigned(202, 8)),
			2332 => std_logic_vector(to_unsigned(58, 8)),
			2333 => std_logic_vector(to_unsigned(156, 8)),
			2334 => std_logic_vector(to_unsigned(33, 8)),
			2335 => std_logic_vector(to_unsigned(117, 8)),
			2336 => std_logic_vector(to_unsigned(18, 8)),
			2337 => std_logic_vector(to_unsigned(213, 8)),
			2338 => std_logic_vector(to_unsigned(68, 8)),
			2339 => std_logic_vector(to_unsigned(215, 8)),
			2340 => std_logic_vector(to_unsigned(50, 8)),
			2341 => std_logic_vector(to_unsigned(217, 8)),
			2342 => std_logic_vector(to_unsigned(175, 8)),
			2343 => std_logic_vector(to_unsigned(82, 8)),
			2344 => std_logic_vector(to_unsigned(1, 8)),
			2345 => std_logic_vector(to_unsigned(181, 8)),
			2346 => std_logic_vector(to_unsigned(161, 8)),
			2347 => std_logic_vector(to_unsigned(34, 8)),
			2348 => std_logic_vector(to_unsigned(123, 8)),
			2349 => std_logic_vector(to_unsigned(63, 8)),
			2350 => std_logic_vector(to_unsigned(114, 8)),
			2351 => std_logic_vector(to_unsigned(19, 8)),
			2352 => std_logic_vector(to_unsigned(163, 8)),
			2353 => std_logic_vector(to_unsigned(188, 8)),
			2354 => std_logic_vector(to_unsigned(52, 8)),
			2355 => std_logic_vector(to_unsigned(95, 8)),
			2356 => std_logic_vector(to_unsigned(74, 8)),
			2357 => std_logic_vector(to_unsigned(28, 8)),
			2358 => std_logic_vector(to_unsigned(52, 8)),
			2359 => std_logic_vector(to_unsigned(250, 8)),
			2360 => std_logic_vector(to_unsigned(109, 8)),
			2361 => std_logic_vector(to_unsigned(82, 8)),
			2362 => std_logic_vector(to_unsigned(48, 8)),
			2363 => std_logic_vector(to_unsigned(103, 8)),
			2364 => std_logic_vector(to_unsigned(179, 8)),
			2365 => std_logic_vector(to_unsigned(50, 8)),
			2366 => std_logic_vector(to_unsigned(217, 8)),
			2367 => std_logic_vector(to_unsigned(65, 8)),
			2368 => std_logic_vector(to_unsigned(247, 8)),
			2369 => std_logic_vector(to_unsigned(174, 8)),
			2370 => std_logic_vector(to_unsigned(189, 8)),
			2371 => std_logic_vector(to_unsigned(62, 8)),
			2372 => std_logic_vector(to_unsigned(122, 8)),
			2373 => std_logic_vector(to_unsigned(45, 8)),
			2374 => std_logic_vector(to_unsigned(238, 8)),
			2375 => std_logic_vector(to_unsigned(91, 8)),
			2376 => std_logic_vector(to_unsigned(177, 8)),
			2377 => std_logic_vector(to_unsigned(186, 8)),
			2378 => std_logic_vector(to_unsigned(240, 8)),
			2379 => std_logic_vector(to_unsigned(178, 8)),
			2380 => std_logic_vector(to_unsigned(76, 8)),
			2381 => std_logic_vector(to_unsigned(98, 8)),
			2382 => std_logic_vector(to_unsigned(153, 8)),
			2383 => std_logic_vector(to_unsigned(112, 8)),
			2384 => std_logic_vector(to_unsigned(251, 8)),
			2385 => std_logic_vector(to_unsigned(243, 8)),
			2386 => std_logic_vector(to_unsigned(76, 8)),
			2387 => std_logic_vector(to_unsigned(102, 8)),
			2388 => std_logic_vector(to_unsigned(70, 8)),
			2389 => std_logic_vector(to_unsigned(102, 8)),
			2390 => std_logic_vector(to_unsigned(56, 8)),
			2391 => std_logic_vector(to_unsigned(214, 8)),
			2392 => std_logic_vector(to_unsigned(111, 8)),
			2393 => std_logic_vector(to_unsigned(88, 8)),
			2394 => std_logic_vector(to_unsigned(50, 8)),
			2395 => std_logic_vector(to_unsigned(205, 8)),
			2396 => std_logic_vector(to_unsigned(146, 8)),
			2397 => std_logic_vector(to_unsigned(210, 8)),
			2398 => std_logic_vector(to_unsigned(206, 8)),
			2399 => std_logic_vector(to_unsigned(97, 8)),
			2400 => std_logic_vector(to_unsigned(197, 8)),
			2401 => std_logic_vector(to_unsigned(181, 8)),
			2402 => std_logic_vector(to_unsigned(167, 8)),
			2403 => std_logic_vector(to_unsigned(107, 8)),
			2404 => std_logic_vector(to_unsigned(114, 8)),
			2405 => std_logic_vector(to_unsigned(230, 8)),
			2406 => std_logic_vector(to_unsigned(44, 8)),
			2407 => std_logic_vector(to_unsigned(70, 8)),
			2408 => std_logic_vector(to_unsigned(190, 8)),
			2409 => std_logic_vector(to_unsigned(173, 8)),
			2410 => std_logic_vector(to_unsigned(180, 8)),
			2411 => std_logic_vector(to_unsigned(148, 8)),
			2412 => std_logic_vector(to_unsigned(130, 8)),
			2413 => std_logic_vector(to_unsigned(112, 8)),
			2414 => std_logic_vector(to_unsigned(90, 8)),
			2415 => std_logic_vector(to_unsigned(40, 8)),
			2416 => std_logic_vector(to_unsigned(36, 8)),
			2417 => std_logic_vector(to_unsigned(141, 8)),
			2418 => std_logic_vector(to_unsigned(55, 8)),
			2419 => std_logic_vector(to_unsigned(196, 8)),
			2420 => std_logic_vector(to_unsigned(166, 8)),
			2421 => std_logic_vector(to_unsigned(20, 8)),
			2422 => std_logic_vector(to_unsigned(209, 8)),
			2423 => std_logic_vector(to_unsigned(141, 8)),
			2424 => std_logic_vector(to_unsigned(21, 8)),
			2425 => std_logic_vector(to_unsigned(206, 8)),
			2426 => std_logic_vector(to_unsigned(28, 8)),
			2427 => std_logic_vector(to_unsigned(209, 8)),
			2428 => std_logic_vector(to_unsigned(184, 8)),
			2429 => std_logic_vector(to_unsigned(102, 8)),
			2430 => std_logic_vector(to_unsigned(191, 8)),
			2431 => std_logic_vector(to_unsigned(155, 8)),
			others => (others => '0'));
component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_rst         : in  std_logic;
      i_start       : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;
begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_rst      	=> tb_rst,
          i_start       => tb_start,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
          o_we 		=> mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;
MEM : process(tb_clk)
begin
    if tb_clk'event and tb_clk = '1' then
        if enable_wire = '1' then
            if mem_we = '1' then
                RAM(conv_integer(mem_address))  <= mem_i_data;
                mem_o_data                      <= mem_i_data after 1 ns;
            else
                mem_o_data <= RAM(conv_integer(mem_address)) after 1 ns;
            end if;
        end if;
    end if;
end process;
test : process is
begin 
    wait for 100 ns;
    wait for c_CLOCK_PERIOD;
    tb_rst <= '1';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_rst <= '0';
    wait for c_CLOCK_PERIOD;
    wait for 100 ns;
    tb_start <= '1';
    wait for c_CLOCK_PERIOD;
    wait until tb_done = '1';
    wait for c_CLOCK_PERIOD;
    tb_start <= '0';
    wait until tb_done = '0';
    wait for 100 ns;
	assert RAM(2432) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(2432))))  severity failure;
	assert RAM(2433) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(2433))))  severity failure;
	assert RAM(2434) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(2434))))  severity failure;
	assert RAM(2435) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(2435))))  severity failure;
	assert RAM(2436) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(2436))))  severity failure;
	assert RAM(2437) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(2437))))  severity failure;
	assert RAM(2438) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(2438))))  severity failure;
	assert RAM(2439) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(2439))))  severity failure;
	assert RAM(2440) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(2440))))  severity failure;
	assert RAM(2441) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(2441))))  severity failure;
	assert RAM(2442) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(2442))))  severity failure;
	assert RAM(2443) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(2443))))  severity failure;
	assert RAM(2444) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(2444))))  severity failure;
	assert RAM(2445) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(2445))))  severity failure;
	assert RAM(2446) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(2446))))  severity failure;
	assert RAM(2447) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(2447))))  severity failure;
	assert RAM(2448) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(2448))))  severity failure;
	assert RAM(2449) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(2449))))  severity failure;
	assert RAM(2450) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(2450))))  severity failure;
	assert RAM(2451) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(2451))))  severity failure;
	assert RAM(2452) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(2452))))  severity failure;
	assert RAM(2453) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(2453))))  severity failure;
	assert RAM(2454) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(2454))))  severity failure;
	assert RAM(2455) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(2455))))  severity failure;
	assert RAM(2456) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(2456))))  severity failure;
	assert RAM(2457) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2457))))  severity failure;
	assert RAM(2458) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(2458))))  severity failure;
	assert RAM(2459) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(2459))))  severity failure;
	assert RAM(2460) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(2460))))  severity failure;
	assert RAM(2461) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2461))))  severity failure;
	assert RAM(2462) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(2462))))  severity failure;
	assert RAM(2463) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(2463))))  severity failure;
	assert RAM(2464) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(2464))))  severity failure;
	assert RAM(2465) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2465))))  severity failure;
	assert RAM(2466) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(2466))))  severity failure;
	assert RAM(2467) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(2467))))  severity failure;
	assert RAM(2468) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2468))))  severity failure;
	assert RAM(2469) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(2469))))  severity failure;
	assert RAM(2470) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(2470))))  severity failure;
	assert RAM(2471) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(2471))))  severity failure;
	assert RAM(2472) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2472))))  severity failure;
	assert RAM(2473) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2473))))  severity failure;
	assert RAM(2474) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(2474))))  severity failure;
	assert RAM(2475) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2475))))  severity failure;
	assert RAM(2476) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(2476))))  severity failure;
	assert RAM(2477) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(2477))))  severity failure;
	assert RAM(2478) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(2478))))  severity failure;
	assert RAM(2479) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2479))))  severity failure;
	assert RAM(2480) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(2480))))  severity failure;
	assert RAM(2481) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(2481))))  severity failure;
	assert RAM(2482) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(2482))))  severity failure;
	assert RAM(2483) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(2483))))  severity failure;
	assert RAM(2484) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(2484))))  severity failure;
	assert RAM(2485) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2485))))  severity failure;
	assert RAM(2486) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(2486))))  severity failure;
	assert RAM(2487) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2487))))  severity failure;
	assert RAM(2488) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(2488))))  severity failure;
	assert RAM(2489) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(2489))))  severity failure;
	assert RAM(2490) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(2490))))  severity failure;
	assert RAM(2491) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(2491))))  severity failure;
	assert RAM(2492) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(2492))))  severity failure;
	assert RAM(2493) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2493))))  severity failure;
	assert RAM(2494) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2494))))  severity failure;
	assert RAM(2495) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(2495))))  severity failure;
	assert RAM(2496) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(2496))))  severity failure;
	assert RAM(2497) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(2497))))  severity failure;
	assert RAM(2498) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(2498))))  severity failure;
	assert RAM(2499) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2499))))  severity failure;
	assert RAM(2500) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(2500))))  severity failure;
	assert RAM(2501) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(2501))))  severity failure;
	assert RAM(2502) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2502))))  severity failure;
	assert RAM(2503) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(2503))))  severity failure;
	assert RAM(2504) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2504))))  severity failure;
	assert RAM(2505) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(2505))))  severity failure;
	assert RAM(2506) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(2506))))  severity failure;
	assert RAM(2507) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(2507))))  severity failure;
	assert RAM(2508) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(2508))))  severity failure;
	assert RAM(2509) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(2509))))  severity failure;
	assert RAM(2510) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(2510))))  severity failure;
	assert RAM(2511) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2511))))  severity failure;
	assert RAM(2512) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2512))))  severity failure;
	assert RAM(2513) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(2513))))  severity failure;
	assert RAM(2514) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(2514))))  severity failure;
	assert RAM(2515) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(2515))))  severity failure;
	assert RAM(2516) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2516))))  severity failure;
	assert RAM(2517) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(2517))))  severity failure;
	assert RAM(2518) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(2518))))  severity failure;
	assert RAM(2519) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(2519))))  severity failure;
	assert RAM(2520) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(2520))))  severity failure;
	assert RAM(2521) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2521))))  severity failure;
	assert RAM(2522) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2522))))  severity failure;
	assert RAM(2523) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(2523))))  severity failure;
	assert RAM(2524) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(2524))))  severity failure;
	assert RAM(2525) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(2525))))  severity failure;
	assert RAM(2526) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(2526))))  severity failure;
	assert RAM(2527) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(2527))))  severity failure;
	assert RAM(2528) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(2528))))  severity failure;
	assert RAM(2529) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(2529))))  severity failure;
	assert RAM(2530) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2530))))  severity failure;
	assert RAM(2531) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(2531))))  severity failure;
	assert RAM(2532) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(2532))))  severity failure;
	assert RAM(2533) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(2533))))  severity failure;
	assert RAM(2534) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(2534))))  severity failure;
	assert RAM(2535) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2535))))  severity failure;
	assert RAM(2536) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2536))))  severity failure;
	assert RAM(2537) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(2537))))  severity failure;
	assert RAM(2538) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2538))))  severity failure;
	assert RAM(2539) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(2539))))  severity failure;
	assert RAM(2540) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(2540))))  severity failure;
	assert RAM(2541) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(2541))))  severity failure;
	assert RAM(2542) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2542))))  severity failure;
	assert RAM(2543) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(2543))))  severity failure;
	assert RAM(2544) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(2544))))  severity failure;
	assert RAM(2545) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(2545))))  severity failure;
	assert RAM(2546) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(2546))))  severity failure;
	assert RAM(2547) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(2547))))  severity failure;
	assert RAM(2548) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2548))))  severity failure;
	assert RAM(2549) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(2549))))  severity failure;
	assert RAM(2550) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2550))))  severity failure;
	assert RAM(2551) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(2551))))  severity failure;
	assert RAM(2552) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2552))))  severity failure;
	assert RAM(2553) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(2553))))  severity failure;
	assert RAM(2554) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(2554))))  severity failure;
	assert RAM(2555) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(2555))))  severity failure;
	assert RAM(2556) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2556))))  severity failure;
	assert RAM(2557) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(2557))))  severity failure;
	assert RAM(2558) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2558))))  severity failure;
	assert RAM(2559) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(2559))))  severity failure;
	assert RAM(2560) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(2560))))  severity failure;
	assert RAM(2561) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(2561))))  severity failure;
	assert RAM(2562) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(2562))))  severity failure;
	assert RAM(2563) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(2563))))  severity failure;
	assert RAM(2564) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(2564))))  severity failure;
	assert RAM(2565) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(2565))))  severity failure;
	assert RAM(2566) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(2566))))  severity failure;
	assert RAM(2567) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(2567))))  severity failure;
	assert RAM(2568) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(2568))))  severity failure;
	assert RAM(2569) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(2569))))  severity failure;
	assert RAM(2570) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2570))))  severity failure;
	assert RAM(2571) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2571))))  severity failure;
	assert RAM(2572) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(2572))))  severity failure;
	assert RAM(2573) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(2573))))  severity failure;
	assert RAM(2574) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2574))))  severity failure;
	assert RAM(2575) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(2575))))  severity failure;
	assert RAM(2576) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(2576))))  severity failure;
	assert RAM(2577) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(2577))))  severity failure;
	assert RAM(2578) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2578))))  severity failure;
	assert RAM(2579) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(2579))))  severity failure;
	assert RAM(2580) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(2580))))  severity failure;
	assert RAM(2581) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(2581))))  severity failure;
	assert RAM(2582) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(2582))))  severity failure;
	assert RAM(2583) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(2583))))  severity failure;
	assert RAM(2584) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(2584))))  severity failure;
	assert RAM(2585) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2585))))  severity failure;
	assert RAM(2586) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2586))))  severity failure;
	assert RAM(2587) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(2587))))  severity failure;
	assert RAM(2588) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(2588))))  severity failure;
	assert RAM(2589) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2589))))  severity failure;
	assert RAM(2590) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(2590))))  severity failure;
	assert RAM(2591) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2591))))  severity failure;
	assert RAM(2592) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(2592))))  severity failure;
	assert RAM(2593) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(2593))))  severity failure;
	assert RAM(2594) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(2594))))  severity failure;
	assert RAM(2595) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(2595))))  severity failure;
	assert RAM(2596) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(2596))))  severity failure;
	assert RAM(2597) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(2597))))  severity failure;
	assert RAM(2598) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2598))))  severity failure;
	assert RAM(2599) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(2599))))  severity failure;
	assert RAM(2600) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(2600))))  severity failure;
	assert RAM(2601) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(2601))))  severity failure;
	assert RAM(2602) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(2602))))  severity failure;
	assert RAM(2603) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(2603))))  severity failure;
	assert RAM(2604) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(2604))))  severity failure;
	assert RAM(2605) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(2605))))  severity failure;
	assert RAM(2606) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(2606))))  severity failure;
	assert RAM(2607) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(2607))))  severity failure;
	assert RAM(2608) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(2608))))  severity failure;
	assert RAM(2609) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2609))))  severity failure;
	assert RAM(2610) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2610))))  severity failure;
	assert RAM(2611) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(2611))))  severity failure;
	assert RAM(2612) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(2612))))  severity failure;
	assert RAM(2613) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(2613))))  severity failure;
	assert RAM(2614) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(2614))))  severity failure;
	assert RAM(2615) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(2615))))  severity failure;
	assert RAM(2616) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2616))))  severity failure;
	assert RAM(2617) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(2617))))  severity failure;
	assert RAM(2618) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(2618))))  severity failure;
	assert RAM(2619) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2619))))  severity failure;
	assert RAM(2620) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(2620))))  severity failure;
	assert RAM(2621) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(2621))))  severity failure;
	assert RAM(2622) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(2622))))  severity failure;
	assert RAM(2623) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(2623))))  severity failure;
	assert RAM(2624) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(2624))))  severity failure;
	assert RAM(2625) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(2625))))  severity failure;
	assert RAM(2626) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(2626))))  severity failure;
	assert RAM(2627) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(2627))))  severity failure;
	assert RAM(2628) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(2628))))  severity failure;
	assert RAM(2629) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(2629))))  severity failure;
	assert RAM(2630) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(2630))))  severity failure;
	assert RAM(2631) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(2631))))  severity failure;
	assert RAM(2632) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(2632))))  severity failure;
	assert RAM(2633) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(2633))))  severity failure;
	assert RAM(2634) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(2634))))  severity failure;
	assert RAM(2635) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(2635))))  severity failure;
	assert RAM(2636) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2636))))  severity failure;
	assert RAM(2637) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(2637))))  severity failure;
	assert RAM(2638) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(2638))))  severity failure;
	assert RAM(2639) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(2639))))  severity failure;
	assert RAM(2640) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2640))))  severity failure;
	assert RAM(2641) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(2641))))  severity failure;
	assert RAM(2642) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(2642))))  severity failure;
	assert RAM(2643) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(2643))))  severity failure;
	assert RAM(2644) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(2644))))  severity failure;
	assert RAM(2645) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(2645))))  severity failure;
	assert RAM(2646) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(2646))))  severity failure;
	assert RAM(2647) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(2647))))  severity failure;
	assert RAM(2648) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2648))))  severity failure;
	assert RAM(2649) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(2649))))  severity failure;
	assert RAM(2650) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(2650))))  severity failure;
	assert RAM(2651) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2651))))  severity failure;
	assert RAM(2652) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(2652))))  severity failure;
	assert RAM(2653) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(2653))))  severity failure;
	assert RAM(2654) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(2654))))  severity failure;
	assert RAM(2655) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(2655))))  severity failure;
	assert RAM(2656) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(2656))))  severity failure;
	assert RAM(2657) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(2657))))  severity failure;
	assert RAM(2658) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(2658))))  severity failure;
	assert RAM(2659) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(2659))))  severity failure;
	assert RAM(2660) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(2660))))  severity failure;
	assert RAM(2661) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(2661))))  severity failure;
	assert RAM(2662) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(2662))))  severity failure;
	assert RAM(2663) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(2663))))  severity failure;
	assert RAM(2664) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(2664))))  severity failure;
	assert RAM(2665) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2665))))  severity failure;
	assert RAM(2666) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(2666))))  severity failure;
	assert RAM(2667) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(2667))))  severity failure;
	assert RAM(2668) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(2668))))  severity failure;
	assert RAM(2669) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(2669))))  severity failure;
	assert RAM(2670) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(2670))))  severity failure;
	assert RAM(2671) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(2671))))  severity failure;
	assert RAM(2672) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(2672))))  severity failure;
	assert RAM(2673) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(2673))))  severity failure;
	assert RAM(2674) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(2674))))  severity failure;
	assert RAM(2675) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(2675))))  severity failure;
	assert RAM(2676) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(2676))))  severity failure;
	assert RAM(2677) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(2677))))  severity failure;
	assert RAM(2678) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(2678))))  severity failure;
	assert RAM(2679) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(2679))))  severity failure;
	assert RAM(2680) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(2680))))  severity failure;
	assert RAM(2681) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(2681))))  severity failure;
	assert RAM(2682) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(2682))))  severity failure;
	assert RAM(2683) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(2683))))  severity failure;
	assert RAM(2684) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(2684))))  severity failure;
	assert RAM(2685) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(2685))))  severity failure;
	assert RAM(2686) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(2686))))  severity failure;
	assert RAM(2687) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(2687))))  severity failure;
	assert RAM(2688) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(2688))))  severity failure;
	assert RAM(2689) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(2689))))  severity failure;
	assert RAM(2690) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2690))))  severity failure;
	assert RAM(2691) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(2691))))  severity failure;
	assert RAM(2692) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(2692))))  severity failure;
	assert RAM(2693) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(2693))))  severity failure;
	assert RAM(2694) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(2694))))  severity failure;
	assert RAM(2695) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(2695))))  severity failure;
	assert RAM(2696) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(2696))))  severity failure;
	assert RAM(2697) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(2697))))  severity failure;
	assert RAM(2698) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(2698))))  severity failure;
	assert RAM(2699) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(2699))))  severity failure;
	assert RAM(2700) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(2700))))  severity failure;
	assert RAM(2701) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(2701))))  severity failure;
	assert RAM(2702) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(2702))))  severity failure;
	assert RAM(2703) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(2703))))  severity failure;
	assert RAM(2704) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2704))))  severity failure;
	assert RAM(2705) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2705))))  severity failure;
	assert RAM(2706) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(2706))))  severity failure;
	assert RAM(2707) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(2707))))  severity failure;
	assert RAM(2708) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(2708))))  severity failure;
	assert RAM(2709) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2709))))  severity failure;
	assert RAM(2710) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2710))))  severity failure;
	assert RAM(2711) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2711))))  severity failure;
	assert RAM(2712) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2712))))  severity failure;
	assert RAM(2713) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(2713))))  severity failure;
	assert RAM(2714) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(2714))))  severity failure;
	assert RAM(2715) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(2715))))  severity failure;
	assert RAM(2716) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(2716))))  severity failure;
	assert RAM(2717) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(2717))))  severity failure;
	assert RAM(2718) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(2718))))  severity failure;
	assert RAM(2719) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2719))))  severity failure;
	assert RAM(2720) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(2720))))  severity failure;
	assert RAM(2721) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(2721))))  severity failure;
	assert RAM(2722) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(2722))))  severity failure;
	assert RAM(2723) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(2723))))  severity failure;
	assert RAM(2724) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(2724))))  severity failure;
	assert RAM(2725) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(2725))))  severity failure;
	assert RAM(2726) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(2726))))  severity failure;
	assert RAM(2727) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(2727))))  severity failure;
	assert RAM(2728) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(2728))))  severity failure;
	assert RAM(2729) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(2729))))  severity failure;
	assert RAM(2730) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(2730))))  severity failure;
	assert RAM(2731) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(2731))))  severity failure;
	assert RAM(2732) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(2732))))  severity failure;
	assert RAM(2733) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(2733))))  severity failure;
	assert RAM(2734) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(2734))))  severity failure;
	assert RAM(2735) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(2735))))  severity failure;
	assert RAM(2736) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(2736))))  severity failure;
	assert RAM(2737) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2737))))  severity failure;
	assert RAM(2738) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(2738))))  severity failure;
	assert RAM(2739) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(2739))))  severity failure;
	assert RAM(2740) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(2740))))  severity failure;
	assert RAM(2741) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(2741))))  severity failure;
	assert RAM(2742) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(2742))))  severity failure;
	assert RAM(2743) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(2743))))  severity failure;
	assert RAM(2744) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(2744))))  severity failure;
	assert RAM(2745) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(2745))))  severity failure;
	assert RAM(2746) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(2746))))  severity failure;
	assert RAM(2747) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(2747))))  severity failure;
	assert RAM(2748) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(2748))))  severity failure;
	assert RAM(2749) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(2749))))  severity failure;
	assert RAM(2750) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(2750))))  severity failure;
	assert RAM(2751) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(2751))))  severity failure;
	assert RAM(2752) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(2752))))  severity failure;
	assert RAM(2753) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2753))))  severity failure;
	assert RAM(2754) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(2754))))  severity failure;
	assert RAM(2755) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(2755))))  severity failure;
	assert RAM(2756) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2756))))  severity failure;
	assert RAM(2757) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(2757))))  severity failure;
	assert RAM(2758) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(2758))))  severity failure;
	assert RAM(2759) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(2759))))  severity failure;
	assert RAM(2760) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2760))))  severity failure;
	assert RAM(2761) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2761))))  severity failure;
	assert RAM(2762) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(2762))))  severity failure;
	assert RAM(2763) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(2763))))  severity failure;
	assert RAM(2764) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(2764))))  severity failure;
	assert RAM(2765) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(2765))))  severity failure;
	assert RAM(2766) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(2766))))  severity failure;
	assert RAM(2767) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(2767))))  severity failure;
	assert RAM(2768) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(2768))))  severity failure;
	assert RAM(2769) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(2769))))  severity failure;
	assert RAM(2770) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(2770))))  severity failure;
	assert RAM(2771) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(2771))))  severity failure;
	assert RAM(2772) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2772))))  severity failure;
	assert RAM(2773) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(2773))))  severity failure;
	assert RAM(2774) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(2774))))  severity failure;
	assert RAM(2775) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(2775))))  severity failure;
	assert RAM(2776) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(2776))))  severity failure;
	assert RAM(2777) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(2777))))  severity failure;
	assert RAM(2778) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(2778))))  severity failure;
	assert RAM(2779) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(2779))))  severity failure;
	assert RAM(2780) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(2780))))  severity failure;
	assert RAM(2781) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(2781))))  severity failure;
	assert RAM(2782) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(2782))))  severity failure;
	assert RAM(2783) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(2783))))  severity failure;
	assert RAM(2784) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2784))))  severity failure;
	assert RAM(2785) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(2785))))  severity failure;
	assert RAM(2786) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(2786))))  severity failure;
	assert RAM(2787) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(2787))))  severity failure;
	assert RAM(2788) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2788))))  severity failure;
	assert RAM(2789) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(2789))))  severity failure;
	assert RAM(2790) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2790))))  severity failure;
	assert RAM(2791) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2791))))  severity failure;
	assert RAM(2792) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(2792))))  severity failure;
	assert RAM(2793) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(2793))))  severity failure;
	assert RAM(2794) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(2794))))  severity failure;
	assert RAM(2795) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2795))))  severity failure;
	assert RAM(2796) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(2796))))  severity failure;
	assert RAM(2797) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(2797))))  severity failure;
	assert RAM(2798) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(2798))))  severity failure;
	assert RAM(2799) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(2799))))  severity failure;
	assert RAM(2800) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(2800))))  severity failure;
	assert RAM(2801) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(2801))))  severity failure;
	assert RAM(2802) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(2802))))  severity failure;
	assert RAM(2803) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(2803))))  severity failure;
	assert RAM(2804) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(2804))))  severity failure;
	assert RAM(2805) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(2805))))  severity failure;
	assert RAM(2806) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(2806))))  severity failure;
	assert RAM(2807) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(2807))))  severity failure;
	assert RAM(2808) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(2808))))  severity failure;
	assert RAM(2809) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(2809))))  severity failure;
	assert RAM(2810) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(2810))))  severity failure;
	assert RAM(2811) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(2811))))  severity failure;
	assert RAM(2812) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(2812))))  severity failure;
	assert RAM(2813) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(2813))))  severity failure;
	assert RAM(2814) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(2814))))  severity failure;
	assert RAM(2815) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(2815))))  severity failure;
	assert RAM(2816) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(2816))))  severity failure;
	assert RAM(2817) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(2817))))  severity failure;
	assert RAM(2818) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(2818))))  severity failure;
	assert RAM(2819) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(2819))))  severity failure;
	assert RAM(2820) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(2820))))  severity failure;
	assert RAM(2821) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(2821))))  severity failure;
	assert RAM(2822) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2822))))  severity failure;
	assert RAM(2823) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(2823))))  severity failure;
	assert RAM(2824) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(2824))))  severity failure;
	assert RAM(2825) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(2825))))  severity failure;
	assert RAM(2826) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(2826))))  severity failure;
	assert RAM(2827) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(2827))))  severity failure;
	assert RAM(2828) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(2828))))  severity failure;
	assert RAM(2829) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(2829))))  severity failure;
	assert RAM(2830) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(2830))))  severity failure;
	assert RAM(2831) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(2831))))  severity failure;
	assert RAM(2832) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(2832))))  severity failure;
	assert RAM(2833) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(2833))))  severity failure;
	assert RAM(2834) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(2834))))  severity failure;
	assert RAM(2835) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(2835))))  severity failure;
	assert RAM(2836) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(2836))))  severity failure;
	assert RAM(2837) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(2837))))  severity failure;
	assert RAM(2838) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(2838))))  severity failure;
	assert RAM(2839) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(2839))))  severity failure;
	assert RAM(2840) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(2840))))  severity failure;
	assert RAM(2841) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(2841))))  severity failure;
	assert RAM(2842) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(2842))))  severity failure;
	assert RAM(2843) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2843))))  severity failure;
	assert RAM(2844) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(2844))))  severity failure;
	assert RAM(2845) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(2845))))  severity failure;
	assert RAM(2846) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(2846))))  severity failure;
	assert RAM(2847) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(2847))))  severity failure;
	assert RAM(2848) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(2848))))  severity failure;
	assert RAM(2849) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2849))))  severity failure;
	assert RAM(2850) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(2850))))  severity failure;
	assert RAM(2851) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(2851))))  severity failure;
	assert RAM(2852) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2852))))  severity failure;
	assert RAM(2853) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(2853))))  severity failure;
	assert RAM(2854) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(2854))))  severity failure;
	assert RAM(2855) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(2855))))  severity failure;
	assert RAM(2856) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(2856))))  severity failure;
	assert RAM(2857) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(2857))))  severity failure;
	assert RAM(2858) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(2858))))  severity failure;
	assert RAM(2859) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(2859))))  severity failure;
	assert RAM(2860) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2860))))  severity failure;
	assert RAM(2861) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(2861))))  severity failure;
	assert RAM(2862) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(2862))))  severity failure;
	assert RAM(2863) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2863))))  severity failure;
	assert RAM(2864) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(2864))))  severity failure;
	assert RAM(2865) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(2865))))  severity failure;
	assert RAM(2866) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2866))))  severity failure;
	assert RAM(2867) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(2867))))  severity failure;
	assert RAM(2868) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(2868))))  severity failure;
	assert RAM(2869) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(2869))))  severity failure;
	assert RAM(2870) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(2870))))  severity failure;
	assert RAM(2871) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(2871))))  severity failure;
	assert RAM(2872) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2872))))  severity failure;
	assert RAM(2873) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(2873))))  severity failure;
	assert RAM(2874) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(2874))))  severity failure;
	assert RAM(2875) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(2875))))  severity failure;
	assert RAM(2876) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(2876))))  severity failure;
	assert RAM(2877) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(2877))))  severity failure;
	assert RAM(2878) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(2878))))  severity failure;
	assert RAM(2879) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2879))))  severity failure;
	assert RAM(2880) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2880))))  severity failure;
	assert RAM(2881) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(2881))))  severity failure;
	assert RAM(2882) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(2882))))  severity failure;
	assert RAM(2883) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2883))))  severity failure;
	assert RAM(2884) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(2884))))  severity failure;
	assert RAM(2885) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(2885))))  severity failure;
	assert RAM(2886) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2886))))  severity failure;
	assert RAM(2887) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(2887))))  severity failure;
	assert RAM(2888) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(2888))))  severity failure;
	assert RAM(2889) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2889))))  severity failure;
	assert RAM(2890) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(2890))))  severity failure;
	assert RAM(2891) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(2891))))  severity failure;
	assert RAM(2892) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(2892))))  severity failure;
	assert RAM(2893) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(2893))))  severity failure;
	assert RAM(2894) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(2894))))  severity failure;
	assert RAM(2895) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(2895))))  severity failure;
	assert RAM(2896) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(2896))))  severity failure;
	assert RAM(2897) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(2897))))  severity failure;
	assert RAM(2898) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(2898))))  severity failure;
	assert RAM(2899) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(2899))))  severity failure;
	assert RAM(2900) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(2900))))  severity failure;
	assert RAM(2901) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(2901))))  severity failure;
	assert RAM(2902) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(2902))))  severity failure;
	assert RAM(2903) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(2903))))  severity failure;
	assert RAM(2904) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(2904))))  severity failure;
	assert RAM(2905) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(2905))))  severity failure;
	assert RAM(2906) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(2906))))  severity failure;
	assert RAM(2907) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(2907))))  severity failure;
	assert RAM(2908) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(2908))))  severity failure;
	assert RAM(2909) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(2909))))  severity failure;
	assert RAM(2910) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(2910))))  severity failure;
	assert RAM(2911) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(2911))))  severity failure;
	assert RAM(2912) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(2912))))  severity failure;
	assert RAM(2913) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(2913))))  severity failure;
	assert RAM(2914) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(2914))))  severity failure;
	assert RAM(2915) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(2915))))  severity failure;
	assert RAM(2916) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(2916))))  severity failure;
	assert RAM(2917) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(2917))))  severity failure;
	assert RAM(2918) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(2918))))  severity failure;
	assert RAM(2919) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(2919))))  severity failure;
	assert RAM(2920) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(2920))))  severity failure;
	assert RAM(2921) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(2921))))  severity failure;
	assert RAM(2922) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(2922))))  severity failure;
	assert RAM(2923) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(2923))))  severity failure;
	assert RAM(2924) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(2924))))  severity failure;
	assert RAM(2925) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(2925))))  severity failure;
	assert RAM(2926) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(2926))))  severity failure;
	assert RAM(2927) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(2927))))  severity failure;
	assert RAM(2928) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(2928))))  severity failure;
	assert RAM(2929) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(2929))))  severity failure;
	assert RAM(2930) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(2930))))  severity failure;
	assert RAM(2931) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2931))))  severity failure;
	assert RAM(2932) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(2932))))  severity failure;
	assert RAM(2933) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(2933))))  severity failure;
	assert RAM(2934) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2934))))  severity failure;
	assert RAM(2935) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(2935))))  severity failure;
	assert RAM(2936) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(2936))))  severity failure;
	assert RAM(2937) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(2937))))  severity failure;
	assert RAM(2938) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(2938))))  severity failure;
	assert RAM(2939) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(2939))))  severity failure;
	assert RAM(2940) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(2940))))  severity failure;
	assert RAM(2941) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2941))))  severity failure;
	assert RAM(2942) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(2942))))  severity failure;
	assert RAM(2943) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2943))))  severity failure;
	assert RAM(2944) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(2944))))  severity failure;
	assert RAM(2945) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(2945))))  severity failure;
	assert RAM(2946) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(2946))))  severity failure;
	assert RAM(2947) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(2947))))  severity failure;
	assert RAM(2948) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(2948))))  severity failure;
	assert RAM(2949) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(2949))))  severity failure;
	assert RAM(2950) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(2950))))  severity failure;
	assert RAM(2951) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(2951))))  severity failure;
	assert RAM(2952) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(2952))))  severity failure;
	assert RAM(2953) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(2953))))  severity failure;
	assert RAM(2954) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(2954))))  severity failure;
	assert RAM(2955) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(2955))))  severity failure;
	assert RAM(2956) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(2956))))  severity failure;
	assert RAM(2957) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(2957))))  severity failure;
	assert RAM(2958) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(2958))))  severity failure;
	assert RAM(2959) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(2959))))  severity failure;
	assert RAM(2960) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(2960))))  severity failure;
	assert RAM(2961) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(2961))))  severity failure;
	assert RAM(2962) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(2962))))  severity failure;
	assert RAM(2963) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(2963))))  severity failure;
	assert RAM(2964) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(2964))))  severity failure;
	assert RAM(2965) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(2965))))  severity failure;
	assert RAM(2966) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(2966))))  severity failure;
	assert RAM(2967) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(2967))))  severity failure;
	assert RAM(2968) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(2968))))  severity failure;
	assert RAM(2969) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(2969))))  severity failure;
	assert RAM(2970) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(2970))))  severity failure;
	assert RAM(2971) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2971))))  severity failure;
	assert RAM(2972) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2972))))  severity failure;
	assert RAM(2973) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(2973))))  severity failure;
	assert RAM(2974) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(2974))))  severity failure;
	assert RAM(2975) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(2975))))  severity failure;
	assert RAM(2976) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(2976))))  severity failure;
	assert RAM(2977) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(2977))))  severity failure;
	assert RAM(2978) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(2978))))  severity failure;
	assert RAM(2979) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(2979))))  severity failure;
	assert RAM(2980) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(2980))))  severity failure;
	assert RAM(2981) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(2981))))  severity failure;
	assert RAM(2982) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(2982))))  severity failure;
	assert RAM(2983) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(2983))))  severity failure;
	assert RAM(2984) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(2984))))  severity failure;
	assert RAM(2985) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(2985))))  severity failure;
	assert RAM(2986) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(2986))))  severity failure;
	assert RAM(2987) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(2987))))  severity failure;
	assert RAM(2988) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(2988))))  severity failure;
	assert RAM(2989) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(2989))))  severity failure;
	assert RAM(2990) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(2990))))  severity failure;
	assert RAM(2991) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(2991))))  severity failure;
	assert RAM(2992) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(2992))))  severity failure;
	assert RAM(2993) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(2993))))  severity failure;
	assert RAM(2994) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(2994))))  severity failure;
	assert RAM(2995) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(2995))))  severity failure;
	assert RAM(2996) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(2996))))  severity failure;
	assert RAM(2997) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(2997))))  severity failure;
	assert RAM(2998) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(2998))))  severity failure;
	assert RAM(2999) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(2999))))  severity failure;
	assert RAM(3000) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(3000))))  severity failure;
	assert RAM(3001) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(3001))))  severity failure;
	assert RAM(3002) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(3002))))  severity failure;
	assert RAM(3003) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(3003))))  severity failure;
	assert RAM(3004) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(3004))))  severity failure;
	assert RAM(3005) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3005))))  severity failure;
	assert RAM(3006) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(3006))))  severity failure;
	assert RAM(3007) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(3007))))  severity failure;
	assert RAM(3008) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(3008))))  severity failure;
	assert RAM(3009) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(3009))))  severity failure;
	assert RAM(3010) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(3010))))  severity failure;
	assert RAM(3011) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(3011))))  severity failure;
	assert RAM(3012) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(3012))))  severity failure;
	assert RAM(3013) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(3013))))  severity failure;
	assert RAM(3014) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(3014))))  severity failure;
	assert RAM(3015) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(3015))))  severity failure;
	assert RAM(3016) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(3016))))  severity failure;
	assert RAM(3017) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(3017))))  severity failure;
	assert RAM(3018) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(3018))))  severity failure;
	assert RAM(3019) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(3019))))  severity failure;
	assert RAM(3020) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3020))))  severity failure;
	assert RAM(3021) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(3021))))  severity failure;
	assert RAM(3022) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(3022))))  severity failure;
	assert RAM(3023) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(3023))))  severity failure;
	assert RAM(3024) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(3024))))  severity failure;
	assert RAM(3025) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(3025))))  severity failure;
	assert RAM(3026) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(3026))))  severity failure;
	assert RAM(3027) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(3027))))  severity failure;
	assert RAM(3028) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(3028))))  severity failure;
	assert RAM(3029) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(3029))))  severity failure;
	assert RAM(3030) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(3030))))  severity failure;
	assert RAM(3031) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(3031))))  severity failure;
	assert RAM(3032) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(3032))))  severity failure;
	assert RAM(3033) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(3033))))  severity failure;
	assert RAM(3034) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(3034))))  severity failure;
	assert RAM(3035) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(3035))))  severity failure;
	assert RAM(3036) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3036))))  severity failure;
	assert RAM(3037) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(3037))))  severity failure;
	assert RAM(3038) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(3038))))  severity failure;
	assert RAM(3039) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(3039))))  severity failure;
	assert RAM(3040) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(3040))))  severity failure;
	assert RAM(3041) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(3041))))  severity failure;
	assert RAM(3042) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(3042))))  severity failure;
	assert RAM(3043) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(3043))))  severity failure;
	assert RAM(3044) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(3044))))  severity failure;
	assert RAM(3045) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(3045))))  severity failure;
	assert RAM(3046) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(3046))))  severity failure;
	assert RAM(3047) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(3047))))  severity failure;
	assert RAM(3048) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(3048))))  severity failure;
	assert RAM(3049) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(3049))))  severity failure;
	assert RAM(3050) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(3050))))  severity failure;
	assert RAM(3051) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(3051))))  severity failure;
	assert RAM(3052) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3052))))  severity failure;
	assert RAM(3053) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(3053))))  severity failure;
	assert RAM(3054) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(3054))))  severity failure;
	assert RAM(3055) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(3055))))  severity failure;
	assert RAM(3056) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(3056))))  severity failure;
	assert RAM(3057) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(3057))))  severity failure;
	assert RAM(3058) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(3058))))  severity failure;
	assert RAM(3059) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(3059))))  severity failure;
	assert RAM(3060) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(3060))))  severity failure;
	assert RAM(3061) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(3061))))  severity failure;
	assert RAM(3062) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3062))))  severity failure;
	assert RAM(3063) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(3063))))  severity failure;
	assert RAM(3064) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(3064))))  severity failure;
	assert RAM(3065) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(3065))))  severity failure;
	assert RAM(3066) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(3066))))  severity failure;
	assert RAM(3067) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(3067))))  severity failure;
	assert RAM(3068) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(3068))))  severity failure;
	assert RAM(3069) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(3069))))  severity failure;
	assert RAM(3070) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(3070))))  severity failure;
	assert RAM(3071) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3071))))  severity failure;
	assert RAM(3072) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(3072))))  severity failure;
	assert RAM(3073) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(3073))))  severity failure;
	assert RAM(3074) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(3074))))  severity failure;
	assert RAM(3075) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3075))))  severity failure;
	assert RAM(3076) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(3076))))  severity failure;
	assert RAM(3077) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(3077))))  severity failure;
	assert RAM(3078) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(3078))))  severity failure;
	assert RAM(3079) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(3079))))  severity failure;
	assert RAM(3080) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(3080))))  severity failure;
	assert RAM(3081) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(3081))))  severity failure;
	assert RAM(3082) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(3082))))  severity failure;
	assert RAM(3083) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(3083))))  severity failure;
	assert RAM(3084) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(3084))))  severity failure;
	assert RAM(3085) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(3085))))  severity failure;
	assert RAM(3086) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(3086))))  severity failure;
	assert RAM(3087) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(3087))))  severity failure;
	assert RAM(3088) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(3088))))  severity failure;
	assert RAM(3089) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(3089))))  severity failure;
	assert RAM(3090) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(3090))))  severity failure;
	assert RAM(3091) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(3091))))  severity failure;
	assert RAM(3092) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(3092))))  severity failure;
	assert RAM(3093) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(3093))))  severity failure;
	assert RAM(3094) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(3094))))  severity failure;
	assert RAM(3095) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(3095))))  severity failure;
	assert RAM(3096) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(3096))))  severity failure;
	assert RAM(3097) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(3097))))  severity failure;
	assert RAM(3098) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(3098))))  severity failure;
	assert RAM(3099) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(3099))))  severity failure;
	assert RAM(3100) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(3100))))  severity failure;
	assert RAM(3101) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(3101))))  severity failure;
	assert RAM(3102) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(3102))))  severity failure;
	assert RAM(3103) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(3103))))  severity failure;
	assert RAM(3104) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(3104))))  severity failure;
	assert RAM(3105) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(3105))))  severity failure;
	assert RAM(3106) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(3106))))  severity failure;
	assert RAM(3107) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(3107))))  severity failure;
	assert RAM(3108) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(3108))))  severity failure;
	assert RAM(3109) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(3109))))  severity failure;
	assert RAM(3110) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(3110))))  severity failure;
	assert RAM(3111) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(3111))))  severity failure;
	assert RAM(3112) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(3112))))  severity failure;
	assert RAM(3113) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(3113))))  severity failure;
	assert RAM(3114) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(3114))))  severity failure;
	assert RAM(3115) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(3115))))  severity failure;
	assert RAM(3116) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(3116))))  severity failure;
	assert RAM(3117) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(3117))))  severity failure;
	assert RAM(3118) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(3118))))  severity failure;
	assert RAM(3119) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(3119))))  severity failure;
	assert RAM(3120) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(3120))))  severity failure;
	assert RAM(3121) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(3121))))  severity failure;
	assert RAM(3122) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(3122))))  severity failure;
	assert RAM(3123) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(3123))))  severity failure;
	assert RAM(3124) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(3124))))  severity failure;
	assert RAM(3125) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(3125))))  severity failure;
	assert RAM(3126) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(3126))))  severity failure;
	assert RAM(3127) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(3127))))  severity failure;
	assert RAM(3128) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(3128))))  severity failure;
	assert RAM(3129) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(3129))))  severity failure;
	assert RAM(3130) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(3130))))  severity failure;
	assert RAM(3131) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(3131))))  severity failure;
	assert RAM(3132) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(3132))))  severity failure;
	assert RAM(3133) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(3133))))  severity failure;
	assert RAM(3134) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(3134))))  severity failure;
	assert RAM(3135) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(3135))))  severity failure;
	assert RAM(3136) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(3136))))  severity failure;
	assert RAM(3137) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(3137))))  severity failure;
	assert RAM(3138) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(3138))))  severity failure;
	assert RAM(3139) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(3139))))  severity failure;
	assert RAM(3140) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(3140))))  severity failure;
	assert RAM(3141) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(3141))))  severity failure;
	assert RAM(3142) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(3142))))  severity failure;
	assert RAM(3143) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(3143))))  severity failure;
	assert RAM(3144) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(3144))))  severity failure;
	assert RAM(3145) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(3145))))  severity failure;
	assert RAM(3146) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(3146))))  severity failure;
	assert RAM(3147) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(3147))))  severity failure;
	assert RAM(3148) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3148))))  severity failure;
	assert RAM(3149) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(3149))))  severity failure;
	assert RAM(3150) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(3150))))  severity failure;
	assert RAM(3151) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(3151))))  severity failure;
	assert RAM(3152) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(3152))))  severity failure;
	assert RAM(3153) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(3153))))  severity failure;
	assert RAM(3154) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(3154))))  severity failure;
	assert RAM(3155) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(3155))))  severity failure;
	assert RAM(3156) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(3156))))  severity failure;
	assert RAM(3157) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(3157))))  severity failure;
	assert RAM(3158) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(3158))))  severity failure;
	assert RAM(3159) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(3159))))  severity failure;
	assert RAM(3160) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(3160))))  severity failure;
	assert RAM(3161) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(3161))))  severity failure;
	assert RAM(3162) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(3162))))  severity failure;
	assert RAM(3163) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(3163))))  severity failure;
	assert RAM(3164) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(3164))))  severity failure;
	assert RAM(3165) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(3165))))  severity failure;
	assert RAM(3166) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(3166))))  severity failure;
	assert RAM(3167) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(3167))))  severity failure;
	assert RAM(3168) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(3168))))  severity failure;
	assert RAM(3169) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3169))))  severity failure;
	assert RAM(3170) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(3170))))  severity failure;
	assert RAM(3171) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(3171))))  severity failure;
	assert RAM(3172) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(3172))))  severity failure;
	assert RAM(3173) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3173))))  severity failure;
	assert RAM(3174) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(3174))))  severity failure;
	assert RAM(3175) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(3175))))  severity failure;
	assert RAM(3176) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(3176))))  severity failure;
	assert RAM(3177) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(3177))))  severity failure;
	assert RAM(3178) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3178))))  severity failure;
	assert RAM(3179) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(3179))))  severity failure;
	assert RAM(3180) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(3180))))  severity failure;
	assert RAM(3181) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(3181))))  severity failure;
	assert RAM(3182) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(3182))))  severity failure;
	assert RAM(3183) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(3183))))  severity failure;
	assert RAM(3184) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(3184))))  severity failure;
	assert RAM(3185) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(3185))))  severity failure;
	assert RAM(3186) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3186))))  severity failure;
	assert RAM(3187) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(3187))))  severity failure;
	assert RAM(3188) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(3188))))  severity failure;
	assert RAM(3189) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(3189))))  severity failure;
	assert RAM(3190) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(3190))))  severity failure;
	assert RAM(3191) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(3191))))  severity failure;
	assert RAM(3192) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(3192))))  severity failure;
	assert RAM(3193) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(3193))))  severity failure;
	assert RAM(3194) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(3194))))  severity failure;
	assert RAM(3195) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(3195))))  severity failure;
	assert RAM(3196) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(3196))))  severity failure;
	assert RAM(3197) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(3197))))  severity failure;
	assert RAM(3198) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(3198))))  severity failure;
	assert RAM(3199) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(3199))))  severity failure;
	assert RAM(3200) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(3200))))  severity failure;
	assert RAM(3201) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(3201))))  severity failure;
	assert RAM(3202) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(3202))))  severity failure;
	assert RAM(3203) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(3203))))  severity failure;
	assert RAM(3204) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(3204))))  severity failure;
	assert RAM(3205) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(3205))))  severity failure;
	assert RAM(3206) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(3206))))  severity failure;
	assert RAM(3207) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(3207))))  severity failure;
	assert RAM(3208) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(3208))))  severity failure;
	assert RAM(3209) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(3209))))  severity failure;
	assert RAM(3210) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(3210))))  severity failure;
	assert RAM(3211) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(3211))))  severity failure;
	assert RAM(3212) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3212))))  severity failure;
	assert RAM(3213) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(3213))))  severity failure;
	assert RAM(3214) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(3214))))  severity failure;
	assert RAM(3215) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(3215))))  severity failure;
	assert RAM(3216) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(3216))))  severity failure;
	assert RAM(3217) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(3217))))  severity failure;
	assert RAM(3218) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(3218))))  severity failure;
	assert RAM(3219) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(3219))))  severity failure;
	assert RAM(3220) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(3220))))  severity failure;
	assert RAM(3221) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(3221))))  severity failure;
	assert RAM(3222) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(3222))))  severity failure;
	assert RAM(3223) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(3223))))  severity failure;
	assert RAM(3224) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(3224))))  severity failure;
	assert RAM(3225) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(3225))))  severity failure;
	assert RAM(3226) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(3226))))  severity failure;
	assert RAM(3227) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(3227))))  severity failure;
	assert RAM(3228) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(3228))))  severity failure;
	assert RAM(3229) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(3229))))  severity failure;
	assert RAM(3230) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(3230))))  severity failure;
	assert RAM(3231) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(3231))))  severity failure;
	assert RAM(3232) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(3232))))  severity failure;
	assert RAM(3233) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(3233))))  severity failure;
	assert RAM(3234) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(3234))))  severity failure;
	assert RAM(3235) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(3235))))  severity failure;
	assert RAM(3236) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(3236))))  severity failure;
	assert RAM(3237) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(3237))))  severity failure;
	assert RAM(3238) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(3238))))  severity failure;
	assert RAM(3239) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(3239))))  severity failure;
	assert RAM(3240) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(3240))))  severity failure;
	assert RAM(3241) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(3241))))  severity failure;
	assert RAM(3242) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(3242))))  severity failure;
	assert RAM(3243) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(3243))))  severity failure;
	assert RAM(3244) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(3244))))  severity failure;
	assert RAM(3245) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(3245))))  severity failure;
	assert RAM(3246) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(3246))))  severity failure;
	assert RAM(3247) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(3247))))  severity failure;
	assert RAM(3248) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(3248))))  severity failure;
	assert RAM(3249) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(3249))))  severity failure;
	assert RAM(3250) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(3250))))  severity failure;
	assert RAM(3251) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(3251))))  severity failure;
	assert RAM(3252) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(3252))))  severity failure;
	assert RAM(3253) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(3253))))  severity failure;
	assert RAM(3254) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(3254))))  severity failure;
	assert RAM(3255) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(3255))))  severity failure;
	assert RAM(3256) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(3256))))  severity failure;
	assert RAM(3257) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(3257))))  severity failure;
	assert RAM(3258) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(3258))))  severity failure;
	assert RAM(3259) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(3259))))  severity failure;
	assert RAM(3260) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(3260))))  severity failure;
	assert RAM(3261) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(3261))))  severity failure;
	assert RAM(3262) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(3262))))  severity failure;
	assert RAM(3263) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(3263))))  severity failure;
	assert RAM(3264) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(3264))))  severity failure;
	assert RAM(3265) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(3265))))  severity failure;
	assert RAM(3266) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(3266))))  severity failure;
	assert RAM(3267) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(3267))))  severity failure;
	assert RAM(3268) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(3268))))  severity failure;
	assert RAM(3269) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(3269))))  severity failure;
	assert RAM(3270) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(3270))))  severity failure;
	assert RAM(3271) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(3271))))  severity failure;
	assert RAM(3272) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(3272))))  severity failure;
	assert RAM(3273) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(3273))))  severity failure;
	assert RAM(3274) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(3274))))  severity failure;
	assert RAM(3275) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(3275))))  severity failure;
	assert RAM(3276) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(3276))))  severity failure;
	assert RAM(3277) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(3277))))  severity failure;
	assert RAM(3278) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(3278))))  severity failure;
	assert RAM(3279) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(3279))))  severity failure;
	assert RAM(3280) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(3280))))  severity failure;
	assert RAM(3281) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(3281))))  severity failure;
	assert RAM(3282) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(3282))))  severity failure;
	assert RAM(3283) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(3283))))  severity failure;
	assert RAM(3284) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(3284))))  severity failure;
	assert RAM(3285) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(3285))))  severity failure;
	assert RAM(3286) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(3286))))  severity failure;
	assert RAM(3287) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(3287))))  severity failure;
	assert RAM(3288) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(3288))))  severity failure;
	assert RAM(3289) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(3289))))  severity failure;
	assert RAM(3290) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(3290))))  severity failure;
	assert RAM(3291) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(3291))))  severity failure;
	assert RAM(3292) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(3292))))  severity failure;
	assert RAM(3293) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(3293))))  severity failure;
	assert RAM(3294) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(3294))))  severity failure;
	assert RAM(3295) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(3295))))  severity failure;
	assert RAM(3296) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(3296))))  severity failure;
	assert RAM(3297) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(3297))))  severity failure;
	assert RAM(3298) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(3298))))  severity failure;
	assert RAM(3299) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(3299))))  severity failure;
	assert RAM(3300) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(3300))))  severity failure;
	assert RAM(3301) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(3301))))  severity failure;
	assert RAM(3302) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(3302))))  severity failure;
	assert RAM(3303) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(3303))))  severity failure;
	assert RAM(3304) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(3304))))  severity failure;
	assert RAM(3305) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(3305))))  severity failure;
	assert RAM(3306) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(3306))))  severity failure;
	assert RAM(3307) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(3307))))  severity failure;
	assert RAM(3308) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(3308))))  severity failure;
	assert RAM(3309) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(3309))))  severity failure;
	assert RAM(3310) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(3310))))  severity failure;
	assert RAM(3311) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(3311))))  severity failure;
	assert RAM(3312) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(3312))))  severity failure;
	assert RAM(3313) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(3313))))  severity failure;
	assert RAM(3314) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(3314))))  severity failure;
	assert RAM(3315) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(3315))))  severity failure;
	assert RAM(3316) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(3316))))  severity failure;
	assert RAM(3317) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(3317))))  severity failure;
	assert RAM(3318) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(3318))))  severity failure;
	assert RAM(3319) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(3319))))  severity failure;
	assert RAM(3320) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(3320))))  severity failure;
	assert RAM(3321) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(3321))))  severity failure;
	assert RAM(3322) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(3322))))  severity failure;
	assert RAM(3323) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(3323))))  severity failure;
	assert RAM(3324) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(3324))))  severity failure;
	assert RAM(3325) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(3325))))  severity failure;
	assert RAM(3326) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(3326))))  severity failure;
	assert RAM(3327) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(3327))))  severity failure;
	assert RAM(3328) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(3328))))  severity failure;
	assert RAM(3329) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(3329))))  severity failure;
	assert RAM(3330) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(3330))))  severity failure;
	assert RAM(3331) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(3331))))  severity failure;
	assert RAM(3332) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(3332))))  severity failure;
	assert RAM(3333) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(3333))))  severity failure;
	assert RAM(3334) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(3334))))  severity failure;
	assert RAM(3335) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(3335))))  severity failure;
	assert RAM(3336) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(3336))))  severity failure;
	assert RAM(3337) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(3337))))  severity failure;
	assert RAM(3338) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(3338))))  severity failure;
	assert RAM(3339) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(3339))))  severity failure;
	assert RAM(3340) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(3340))))  severity failure;
	assert RAM(3341) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(3341))))  severity failure;
	assert RAM(3342) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(3342))))  severity failure;
	assert RAM(3343) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(3343))))  severity failure;
	assert RAM(3344) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(3344))))  severity failure;
	assert RAM(3345) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3345))))  severity failure;
	assert RAM(3346) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(3346))))  severity failure;
	assert RAM(3347) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(3347))))  severity failure;
	assert RAM(3348) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(3348))))  severity failure;
	assert RAM(3349) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(3349))))  severity failure;
	assert RAM(3350) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(3350))))  severity failure;
	assert RAM(3351) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(3351))))  severity failure;
	assert RAM(3352) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(3352))))  severity failure;
	assert RAM(3353) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(3353))))  severity failure;
	assert RAM(3354) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(3354))))  severity failure;
	assert RAM(3355) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(3355))))  severity failure;
	assert RAM(3356) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(3356))))  severity failure;
	assert RAM(3357) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(3357))))  severity failure;
	assert RAM(3358) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(3358))))  severity failure;
	assert RAM(3359) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(3359))))  severity failure;
	assert RAM(3360) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(3360))))  severity failure;
	assert RAM(3361) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(3361))))  severity failure;
	assert RAM(3362) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3362))))  severity failure;
	assert RAM(3363) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3363))))  severity failure;
	assert RAM(3364) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(3364))))  severity failure;
	assert RAM(3365) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(3365))))  severity failure;
	assert RAM(3366) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3366))))  severity failure;
	assert RAM(3367) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(3367))))  severity failure;
	assert RAM(3368) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(3368))))  severity failure;
	assert RAM(3369) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(3369))))  severity failure;
	assert RAM(3370) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(3370))))  severity failure;
	assert RAM(3371) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(3371))))  severity failure;
	assert RAM(3372) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(3372))))  severity failure;
	assert RAM(3373) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(3373))))  severity failure;
	assert RAM(3374) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(3374))))  severity failure;
	assert RAM(3375) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(3375))))  severity failure;
	assert RAM(3376) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(3376))))  severity failure;
	assert RAM(3377) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(3377))))  severity failure;
	assert RAM(3378) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3378))))  severity failure;
	assert RAM(3379) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(3379))))  severity failure;
	assert RAM(3380) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(3380))))  severity failure;
	assert RAM(3381) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(3381))))  severity failure;
	assert RAM(3382) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(3382))))  severity failure;
	assert RAM(3383) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(3383))))  severity failure;
	assert RAM(3384) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(3384))))  severity failure;
	assert RAM(3385) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(3385))))  severity failure;
	assert RAM(3386) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(3386))))  severity failure;
	assert RAM(3387) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(3387))))  severity failure;
	assert RAM(3388) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(3388))))  severity failure;
	assert RAM(3389) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(3389))))  severity failure;
	assert RAM(3390) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(3390))))  severity failure;
	assert RAM(3391) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(3391))))  severity failure;
	assert RAM(3392) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(3392))))  severity failure;
	assert RAM(3393) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(3393))))  severity failure;
	assert RAM(3394) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(3394))))  severity failure;
	assert RAM(3395) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(3395))))  severity failure;
	assert RAM(3396) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(3396))))  severity failure;
	assert RAM(3397) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(3397))))  severity failure;
	assert RAM(3398) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(3398))))  severity failure;
	assert RAM(3399) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(3399))))  severity failure;
	assert RAM(3400) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(3400))))  severity failure;
	assert RAM(3401) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(3401))))  severity failure;
	assert RAM(3402) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(3402))))  severity failure;
	assert RAM(3403) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(3403))))  severity failure;
	assert RAM(3404) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(3404))))  severity failure;
	assert RAM(3405) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(3405))))  severity failure;
	assert RAM(3406) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(3406))))  severity failure;
	assert RAM(3407) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(3407))))  severity failure;
	assert RAM(3408) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(3408))))  severity failure;
	assert RAM(3409) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(3409))))  severity failure;
	assert RAM(3410) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3410))))  severity failure;
	assert RAM(3411) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(3411))))  severity failure;
	assert RAM(3412) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(3412))))  severity failure;
	assert RAM(3413) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(3413))))  severity failure;
	assert RAM(3414) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(3414))))  severity failure;
	assert RAM(3415) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(3415))))  severity failure;
	assert RAM(3416) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(3416))))  severity failure;
	assert RAM(3417) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(3417))))  severity failure;
	assert RAM(3418) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(3418))))  severity failure;
	assert RAM(3419) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(3419))))  severity failure;
	assert RAM(3420) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(3420))))  severity failure;
	assert RAM(3421) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(3421))))  severity failure;
	assert RAM(3422) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(3422))))  severity failure;
	assert RAM(3423) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(3423))))  severity failure;
	assert RAM(3424) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(3424))))  severity failure;
	assert RAM(3425) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(3425))))  severity failure;
	assert RAM(3426) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(3426))))  severity failure;
	assert RAM(3427) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(3427))))  severity failure;
	assert RAM(3428) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(3428))))  severity failure;
	assert RAM(3429) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(3429))))  severity failure;
	assert RAM(3430) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(3430))))  severity failure;
	assert RAM(3431) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(3431))))  severity failure;
	assert RAM(3432) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(3432))))  severity failure;
	assert RAM(3433) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(3433))))  severity failure;
	assert RAM(3434) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(3434))))  severity failure;
	assert RAM(3435) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(3435))))  severity failure;
	assert RAM(3436) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(3436))))  severity failure;
	assert RAM(3437) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(3437))))  severity failure;
	assert RAM(3438) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(3438))))  severity failure;
	assert RAM(3439) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(3439))))  severity failure;
	assert RAM(3440) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(3440))))  severity failure;
	assert RAM(3441) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(3441))))  severity failure;
	assert RAM(3442) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(3442))))  severity failure;
	assert RAM(3443) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(3443))))  severity failure;
	assert RAM(3444) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(3444))))  severity failure;
	assert RAM(3445) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(3445))))  severity failure;
	assert RAM(3446) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(3446))))  severity failure;
	assert RAM(3447) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(3447))))  severity failure;
	assert RAM(3448) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(3448))))  severity failure;
	assert RAM(3449) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(3449))))  severity failure;
	assert RAM(3450) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(3450))))  severity failure;
	assert RAM(3451) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(3451))))  severity failure;
	assert RAM(3452) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(3452))))  severity failure;
	assert RAM(3453) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(3453))))  severity failure;
	assert RAM(3454) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(3454))))  severity failure;
	assert RAM(3455) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(3455))))  severity failure;
	assert RAM(3456) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(3456))))  severity failure;
	assert RAM(3457) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(3457))))  severity failure;
	assert RAM(3458) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(3458))))  severity failure;
	assert RAM(3459) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(3459))))  severity failure;
	assert RAM(3460) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(3460))))  severity failure;
	assert RAM(3461) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(3461))))  severity failure;
	assert RAM(3462) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(3462))))  severity failure;
	assert RAM(3463) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(3463))))  severity failure;
	assert RAM(3464) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(3464))))  severity failure;
	assert RAM(3465) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(3465))))  severity failure;
	assert RAM(3466) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3466))))  severity failure;
	assert RAM(3467) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(3467))))  severity failure;
	assert RAM(3468) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(3468))))  severity failure;
	assert RAM(3469) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(3469))))  severity failure;
	assert RAM(3470) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(3470))))  severity failure;
	assert RAM(3471) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3471))))  severity failure;
	assert RAM(3472) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(3472))))  severity failure;
	assert RAM(3473) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3473))))  severity failure;
	assert RAM(3474) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(3474))))  severity failure;
	assert RAM(3475) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(3475))))  severity failure;
	assert RAM(3476) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(3476))))  severity failure;
	assert RAM(3477) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(3477))))  severity failure;
	assert RAM(3478) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(3478))))  severity failure;
	assert RAM(3479) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(3479))))  severity failure;
	assert RAM(3480) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(3480))))  severity failure;
	assert RAM(3481) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(3481))))  severity failure;
	assert RAM(3482) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(3482))))  severity failure;
	assert RAM(3483) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(3483))))  severity failure;
	assert RAM(3484) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(3484))))  severity failure;
	assert RAM(3485) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(3485))))  severity failure;
	assert RAM(3486) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(3486))))  severity failure;
	assert RAM(3487) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(3487))))  severity failure;
	assert RAM(3488) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(3488))))  severity failure;
	assert RAM(3489) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(3489))))  severity failure;
	assert RAM(3490) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3490))))  severity failure;
	assert RAM(3491) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(3491))))  severity failure;
	assert RAM(3492) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(3492))))  severity failure;
	assert RAM(3493) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(3493))))  severity failure;
	assert RAM(3494) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(3494))))  severity failure;
	assert RAM(3495) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(3495))))  severity failure;
	assert RAM(3496) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(3496))))  severity failure;
	assert RAM(3497) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3497))))  severity failure;
	assert RAM(3498) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(3498))))  severity failure;
	assert RAM(3499) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(3499))))  severity failure;
	assert RAM(3500) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(3500))))  severity failure;
	assert RAM(3501) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(3501))))  severity failure;
	assert RAM(3502) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(3502))))  severity failure;
	assert RAM(3503) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3503))))  severity failure;
	assert RAM(3504) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(3504))))  severity failure;
	assert RAM(3505) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(3505))))  severity failure;
	assert RAM(3506) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(3506))))  severity failure;
	assert RAM(3507) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(3507))))  severity failure;
	assert RAM(3508) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(3508))))  severity failure;
	assert RAM(3509) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(3509))))  severity failure;
	assert RAM(3510) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(3510))))  severity failure;
	assert RAM(3511) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(3511))))  severity failure;
	assert RAM(3512) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(3512))))  severity failure;
	assert RAM(3513) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(3513))))  severity failure;
	assert RAM(3514) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(3514))))  severity failure;
	assert RAM(3515) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(3515))))  severity failure;
	assert RAM(3516) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(3516))))  severity failure;
	assert RAM(3517) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(3517))))  severity failure;
	assert RAM(3518) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(3518))))  severity failure;
	assert RAM(3519) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(3519))))  severity failure;
	assert RAM(3520) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(3520))))  severity failure;
	assert RAM(3521) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(3521))))  severity failure;
	assert RAM(3522) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(3522))))  severity failure;
	assert RAM(3523) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(3523))))  severity failure;
	assert RAM(3524) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(3524))))  severity failure;
	assert RAM(3525) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(3525))))  severity failure;
	assert RAM(3526) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(3526))))  severity failure;
	assert RAM(3527) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(3527))))  severity failure;
	assert RAM(3528) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(3528))))  severity failure;
	assert RAM(3529) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(3529))))  severity failure;
	assert RAM(3530) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(3530))))  severity failure;
	assert RAM(3531) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(3531))))  severity failure;
	assert RAM(3532) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(3532))))  severity failure;
	assert RAM(3533) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(3533))))  severity failure;
	assert RAM(3534) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(3534))))  severity failure;
	assert RAM(3535) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(3535))))  severity failure;
	assert RAM(3536) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(3536))))  severity failure;
	assert RAM(3537) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(3537))))  severity failure;
	assert RAM(3538) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(3538))))  severity failure;
	assert RAM(3539) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(3539))))  severity failure;
	assert RAM(3540) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(3540))))  severity failure;
	assert RAM(3541) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(3541))))  severity failure;
	assert RAM(3542) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(3542))))  severity failure;
	assert RAM(3543) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(3543))))  severity failure;
	assert RAM(3544) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(3544))))  severity failure;
	assert RAM(3545) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(3545))))  severity failure;
	assert RAM(3546) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(3546))))  severity failure;
	assert RAM(3547) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(3547))))  severity failure;
	assert RAM(3548) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(3548))))  severity failure;
	assert RAM(3549) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(3549))))  severity failure;
	assert RAM(3550) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(3550))))  severity failure;
	assert RAM(3551) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3551))))  severity failure;
	assert RAM(3552) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(3552))))  severity failure;
	assert RAM(3553) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(3553))))  severity failure;
	assert RAM(3554) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3554))))  severity failure;
	assert RAM(3555) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(3555))))  severity failure;
	assert RAM(3556) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(3556))))  severity failure;
	assert RAM(3557) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(3557))))  severity failure;
	assert RAM(3558) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(3558))))  severity failure;
	assert RAM(3559) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(3559))))  severity failure;
	assert RAM(3560) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(3560))))  severity failure;
	assert RAM(3561) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(3561))))  severity failure;
	assert RAM(3562) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(3562))))  severity failure;
	assert RAM(3563) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(3563))))  severity failure;
	assert RAM(3564) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(3564))))  severity failure;
	assert RAM(3565) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(3565))))  severity failure;
	assert RAM(3566) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(3566))))  severity failure;
	assert RAM(3567) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(3567))))  severity failure;
	assert RAM(3568) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(3568))))  severity failure;
	assert RAM(3569) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(3569))))  severity failure;
	assert RAM(3570) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(3570))))  severity failure;
	assert RAM(3571) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(3571))))  severity failure;
	assert RAM(3572) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(3572))))  severity failure;
	assert RAM(3573) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(3573))))  severity failure;
	assert RAM(3574) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(3574))))  severity failure;
	assert RAM(3575) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(3575))))  severity failure;
	assert RAM(3576) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(3576))))  severity failure;
	assert RAM(3577) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(3577))))  severity failure;
	assert RAM(3578) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(3578))))  severity failure;
	assert RAM(3579) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(3579))))  severity failure;
	assert RAM(3580) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(3580))))  severity failure;
	assert RAM(3581) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(3581))))  severity failure;
	assert RAM(3582) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(3582))))  severity failure;
	assert RAM(3583) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(3583))))  severity failure;
	assert RAM(3584) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(3584))))  severity failure;
	assert RAM(3585) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(3585))))  severity failure;
	assert RAM(3586) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(3586))))  severity failure;
	assert RAM(3587) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(3587))))  severity failure;
	assert RAM(3588) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(3588))))  severity failure;
	assert RAM(3589) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(3589))))  severity failure;
	assert RAM(3590) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(3590))))  severity failure;
	assert RAM(3591) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(3591))))  severity failure;
	assert RAM(3592) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(3592))))  severity failure;
	assert RAM(3593) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(3593))))  severity failure;
	assert RAM(3594) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(3594))))  severity failure;
	assert RAM(3595) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(3595))))  severity failure;
	assert RAM(3596) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(3596))))  severity failure;
	assert RAM(3597) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(3597))))  severity failure;
	assert RAM(3598) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(3598))))  severity failure;
	assert RAM(3599) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(3599))))  severity failure;
	assert RAM(3600) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(3600))))  severity failure;
	assert RAM(3601) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(3601))))  severity failure;
	assert RAM(3602) = std_logic_vector(to_unsigned(51, 8)) report "TEST FALLITO (WORKING ZONE). Expected  51  found " & integer'image(to_integer(unsigned(RAM(3602))))  severity failure;
	assert RAM(3603) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(3603))))  severity failure;
	assert RAM(3604) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(3604))))  severity failure;
	assert RAM(3605) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(3605))))  severity failure;
	assert RAM(3606) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(3606))))  severity failure;
	assert RAM(3607) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(3607))))  severity failure;
	assert RAM(3608) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(3608))))  severity failure;
	assert RAM(3609) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(3609))))  severity failure;
	assert RAM(3610) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(3610))))  severity failure;
	assert RAM(3611) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(3611))))  severity failure;
	assert RAM(3612) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(3612))))  severity failure;
	assert RAM(3613) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(3613))))  severity failure;
	assert RAM(3614) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(3614))))  severity failure;
	assert RAM(3615) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(3615))))  severity failure;
	assert RAM(3616) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(3616))))  severity failure;
	assert RAM(3617) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(3617))))  severity failure;
	assert RAM(3618) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(3618))))  severity failure;
	assert RAM(3619) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(3619))))  severity failure;
	assert RAM(3620) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(3620))))  severity failure;
	assert RAM(3621) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(3621))))  severity failure;
	assert RAM(3622) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(3622))))  severity failure;
	assert RAM(3623) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(3623))))  severity failure;
	assert RAM(3624) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(3624))))  severity failure;
	assert RAM(3625) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(3625))))  severity failure;
	assert RAM(3626) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(3626))))  severity failure;
	assert RAM(3627) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(3627))))  severity failure;
	assert RAM(3628) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(3628))))  severity failure;
	assert RAM(3629) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(3629))))  severity failure;
	assert RAM(3630) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(3630))))  severity failure;
	assert RAM(3631) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(3631))))  severity failure;
	assert RAM(3632) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(3632))))  severity failure;
	assert RAM(3633) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(3633))))  severity failure;
	assert RAM(3634) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(3634))))  severity failure;
	assert RAM(3635) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(3635))))  severity failure;
	assert RAM(3636) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(3636))))  severity failure;
	assert RAM(3637) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(3637))))  severity failure;
	assert RAM(3638) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(3638))))  severity failure;
	assert RAM(3639) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(3639))))  severity failure;
	assert RAM(3640) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(3640))))  severity failure;
	assert RAM(3641) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(3641))))  severity failure;
	assert RAM(3642) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(3642))))  severity failure;
	assert RAM(3643) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(3643))))  severity failure;
	assert RAM(3644) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(3644))))  severity failure;
	assert RAM(3645) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(3645))))  severity failure;
	assert RAM(3646) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(3646))))  severity failure;
	assert RAM(3647) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(3647))))  severity failure;
	assert RAM(3648) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(3648))))  severity failure;
	assert RAM(3649) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(3649))))  severity failure;
	assert RAM(3650) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(3650))))  severity failure;
	assert RAM(3651) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(3651))))  severity failure;
	assert RAM(3652) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3652))))  severity failure;
	assert RAM(3653) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(3653))))  severity failure;
	assert RAM(3654) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(3654))))  severity failure;
	assert RAM(3655) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(3655))))  severity failure;
	assert RAM(3656) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(3656))))  severity failure;
	assert RAM(3657) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(3657))))  severity failure;
	assert RAM(3658) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(3658))))  severity failure;
	assert RAM(3659) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(3659))))  severity failure;
	assert RAM(3660) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(3660))))  severity failure;
	assert RAM(3661) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(3661))))  severity failure;
	assert RAM(3662) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(3662))))  severity failure;
	assert RAM(3663) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(3663))))  severity failure;
	assert RAM(3664) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(3664))))  severity failure;
	assert RAM(3665) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(3665))))  severity failure;
	assert RAM(3666) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3666))))  severity failure;
	assert RAM(3667) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(3667))))  severity failure;
	assert RAM(3668) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(3668))))  severity failure;
	assert RAM(3669) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(3669))))  severity failure;
	assert RAM(3670) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(3670))))  severity failure;
	assert RAM(3671) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(3671))))  severity failure;
	assert RAM(3672) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(3672))))  severity failure;
	assert RAM(3673) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(3673))))  severity failure;
	assert RAM(3674) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(3674))))  severity failure;
	assert RAM(3675) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(3675))))  severity failure;
	assert RAM(3676) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(3676))))  severity failure;
	assert RAM(3677) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(3677))))  severity failure;
	assert RAM(3678) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(3678))))  severity failure;
	assert RAM(3679) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(3679))))  severity failure;
	assert RAM(3680) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(3680))))  severity failure;
	assert RAM(3681) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(3681))))  severity failure;
	assert RAM(3682) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(3682))))  severity failure;
	assert RAM(3683) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(3683))))  severity failure;
	assert RAM(3684) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(3684))))  severity failure;
	assert RAM(3685) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(3685))))  severity failure;
	assert RAM(3686) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(3686))))  severity failure;
	assert RAM(3687) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(3687))))  severity failure;
	assert RAM(3688) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(3688))))  severity failure;
	assert RAM(3689) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(3689))))  severity failure;
	assert RAM(3690) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(3690))))  severity failure;
	assert RAM(3691) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(3691))))  severity failure;
	assert RAM(3692) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(3692))))  severity failure;
	assert RAM(3693) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(3693))))  severity failure;
	assert RAM(3694) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(3694))))  severity failure;
	assert RAM(3695) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3695))))  severity failure;
	assert RAM(3696) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(3696))))  severity failure;
	assert RAM(3697) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(3697))))  severity failure;
	assert RAM(3698) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(3698))))  severity failure;
	assert RAM(3699) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(3699))))  severity failure;
	assert RAM(3700) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(3700))))  severity failure;
	assert RAM(3701) = std_logic_vector(to_unsigned(8, 8)) report "TEST FALLITO (WORKING ZONE). Expected  8  found " & integer'image(to_integer(unsigned(RAM(3701))))  severity failure;
	assert RAM(3702) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(3702))))  severity failure;
	assert RAM(3703) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(3703))))  severity failure;
	assert RAM(3704) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3704))))  severity failure;
	assert RAM(3705) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(3705))))  severity failure;
	assert RAM(3706) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(3706))))  severity failure;
	assert RAM(3707) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3707))))  severity failure;
	assert RAM(3708) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(3708))))  severity failure;
	assert RAM(3709) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(3709))))  severity failure;
	assert RAM(3710) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(3710))))  severity failure;
	assert RAM(3711) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(3711))))  severity failure;
	assert RAM(3712) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(3712))))  severity failure;
	assert RAM(3713) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(3713))))  severity failure;
	assert RAM(3714) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(3714))))  severity failure;
	assert RAM(3715) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(3715))))  severity failure;
	assert RAM(3716) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(3716))))  severity failure;
	assert RAM(3717) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(3717))))  severity failure;
	assert RAM(3718) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(3718))))  severity failure;
	assert RAM(3719) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(3719))))  severity failure;
	assert RAM(3720) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(3720))))  severity failure;
	assert RAM(3721) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(3721))))  severity failure;
	assert RAM(3722) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(3722))))  severity failure;
	assert RAM(3723) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(3723))))  severity failure;
	assert RAM(3724) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(3724))))  severity failure;
	assert RAM(3725) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(3725))))  severity failure;
	assert RAM(3726) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(3726))))  severity failure;
	assert RAM(3727) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(3727))))  severity failure;
	assert RAM(3728) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(3728))))  severity failure;
	assert RAM(3729) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(3729))))  severity failure;
	assert RAM(3730) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(3730))))  severity failure;
	assert RAM(3731) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(3731))))  severity failure;
	assert RAM(3732) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(3732))))  severity failure;
	assert RAM(3733) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(3733))))  severity failure;
	assert RAM(3734) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(3734))))  severity failure;
	assert RAM(3735) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(3735))))  severity failure;
	assert RAM(3736) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(3736))))  severity failure;
	assert RAM(3737) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(3737))))  severity failure;
	assert RAM(3738) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(3738))))  severity failure;
	assert RAM(3739) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3739))))  severity failure;
	assert RAM(3740) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(3740))))  severity failure;
	assert RAM(3741) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(3741))))  severity failure;
	assert RAM(3742) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(3742))))  severity failure;
	assert RAM(3743) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(3743))))  severity failure;
	assert RAM(3744) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(3744))))  severity failure;
	assert RAM(3745) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(3745))))  severity failure;
	assert RAM(3746) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(3746))))  severity failure;
	assert RAM(3747) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(3747))))  severity failure;
	assert RAM(3748) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3748))))  severity failure;
	assert RAM(3749) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(3749))))  severity failure;
	assert RAM(3750) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(3750))))  severity failure;
	assert RAM(3751) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(3751))))  severity failure;
	assert RAM(3752) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(3752))))  severity failure;
	assert RAM(3753) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(3753))))  severity failure;
	assert RAM(3754) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(3754))))  severity failure;
	assert RAM(3755) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(3755))))  severity failure;
	assert RAM(3756) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(3756))))  severity failure;
	assert RAM(3757) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(3757))))  severity failure;
	assert RAM(3758) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(3758))))  severity failure;
	assert RAM(3759) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3759))))  severity failure;
	assert RAM(3760) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(3760))))  severity failure;
	assert RAM(3761) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(3761))))  severity failure;
	assert RAM(3762) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3762))))  severity failure;
	assert RAM(3763) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(3763))))  severity failure;
	assert RAM(3764) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(3764))))  severity failure;
	assert RAM(3765) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(3765))))  severity failure;
	assert RAM(3766) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(3766))))  severity failure;
	assert RAM(3767) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(3767))))  severity failure;
	assert RAM(3768) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(3768))))  severity failure;
	assert RAM(3769) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3769))))  severity failure;
	assert RAM(3770) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(3770))))  severity failure;
	assert RAM(3771) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(3771))))  severity failure;
	assert RAM(3772) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(3772))))  severity failure;
	assert RAM(3773) = std_logic_vector(to_unsigned(77, 8)) report "TEST FALLITO (WORKING ZONE). Expected  77  found " & integer'image(to_integer(unsigned(RAM(3773))))  severity failure;
	assert RAM(3774) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(3774))))  severity failure;
	assert RAM(3775) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(3775))))  severity failure;
	assert RAM(3776) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(3776))))  severity failure;
	assert RAM(3777) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(3777))))  severity failure;
	assert RAM(3778) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(3778))))  severity failure;
	assert RAM(3779) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(3779))))  severity failure;
	assert RAM(3780) = std_logic_vector(to_unsigned(43, 8)) report "TEST FALLITO (WORKING ZONE). Expected  43  found " & integer'image(to_integer(unsigned(RAM(3780))))  severity failure;
	assert RAM(3781) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(3781))))  severity failure;
	assert RAM(3782) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(3782))))  severity failure;
	assert RAM(3783) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(3783))))  severity failure;
	assert RAM(3784) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(3784))))  severity failure;
	assert RAM(3785) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(3785))))  severity failure;
	assert RAM(3786) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(3786))))  severity failure;
	assert RAM(3787) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(3787))))  severity failure;
	assert RAM(3788) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(3788))))  severity failure;
	assert RAM(3789) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(3789))))  severity failure;
	assert RAM(3790) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(3790))))  severity failure;
	assert RAM(3791) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(3791))))  severity failure;
	assert RAM(3792) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(3792))))  severity failure;
	assert RAM(3793) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(3793))))  severity failure;
	assert RAM(3794) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(3794))))  severity failure;
	assert RAM(3795) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(3795))))  severity failure;
	assert RAM(3796) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(3796))))  severity failure;
	assert RAM(3797) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(3797))))  severity failure;
	assert RAM(3798) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(3798))))  severity failure;
	assert RAM(3799) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(3799))))  severity failure;
	assert RAM(3800) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(3800))))  severity failure;
	assert RAM(3801) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(3801))))  severity failure;
	assert RAM(3802) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(3802))))  severity failure;
	assert RAM(3803) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(3803))))  severity failure;
	assert RAM(3804) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(3804))))  severity failure;
	assert RAM(3805) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(3805))))  severity failure;
	assert RAM(3806) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(3806))))  severity failure;
	assert RAM(3807) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(3807))))  severity failure;
	assert RAM(3808) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(3808))))  severity failure;
	assert RAM(3809) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(3809))))  severity failure;
	assert RAM(3810) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(3810))))  severity failure;
	assert RAM(3811) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(3811))))  severity failure;
	assert RAM(3812) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(3812))))  severity failure;
	assert RAM(3813) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(3813))))  severity failure;
	assert RAM(3814) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(3814))))  severity failure;
	assert RAM(3815) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(3815))))  severity failure;
	assert RAM(3816) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(3816))))  severity failure;
	assert RAM(3817) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(3817))))  severity failure;
	assert RAM(3818) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(3818))))  severity failure;
	assert RAM(3819) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(3819))))  severity failure;
	assert RAM(3820) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(3820))))  severity failure;
	assert RAM(3821) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(3821))))  severity failure;
	assert RAM(3822) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(3822))))  severity failure;
	assert RAM(3823) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(3823))))  severity failure;
	assert RAM(3824) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(3824))))  severity failure;
	assert RAM(3825) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(3825))))  severity failure;
	assert RAM(3826) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(3826))))  severity failure;
	assert RAM(3827) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(3827))))  severity failure;
	assert RAM(3828) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(3828))))  severity failure;
	assert RAM(3829) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(3829))))  severity failure;
	assert RAM(3830) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(3830))))  severity failure;
	assert RAM(3831) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(3831))))  severity failure;
	assert RAM(3832) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(3832))))  severity failure;
	assert RAM(3833) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(3833))))  severity failure;
	assert RAM(3834) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(3834))))  severity failure;
	assert RAM(3835) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(3835))))  severity failure;
	assert RAM(3836) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(3836))))  severity failure;
	assert RAM(3837) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(3837))))  severity failure;
	assert RAM(3838) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(3838))))  severity failure;
	assert RAM(3839) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(3839))))  severity failure;
	assert RAM(3840) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(3840))))  severity failure;
	assert RAM(3841) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(3841))))  severity failure;
	assert RAM(3842) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(3842))))  severity failure;
	assert RAM(3843) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(3843))))  severity failure;
	assert RAM(3844) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(3844))))  severity failure;
	assert RAM(3845) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(3845))))  severity failure;
	assert RAM(3846) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(3846))))  severity failure;
	assert RAM(3847) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(3847))))  severity failure;
	assert RAM(3848) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(3848))))  severity failure;
	assert RAM(3849) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(3849))))  severity failure;
	assert RAM(3850) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(3850))))  severity failure;
	assert RAM(3851) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(3851))))  severity failure;
	assert RAM(3852) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(3852))))  severity failure;
	assert RAM(3853) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(3853))))  severity failure;
	assert RAM(3854) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(3854))))  severity failure;
	assert RAM(3855) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(3855))))  severity failure;
	assert RAM(3856) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(3856))))  severity failure;
	assert RAM(3857) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(3857))))  severity failure;
	assert RAM(3858) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(3858))))  severity failure;
	assert RAM(3859) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(3859))))  severity failure;
	assert RAM(3860) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(3860))))  severity failure;
	assert RAM(3861) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(3861))))  severity failure;
	assert RAM(3862) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(3862))))  severity failure;
	assert RAM(3863) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(3863))))  severity failure;
	assert RAM(3864) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(3864))))  severity failure;
	assert RAM(3865) = std_logic_vector(to_unsigned(176, 8)) report "TEST FALLITO (WORKING ZONE). Expected  176  found " & integer'image(to_integer(unsigned(RAM(3865))))  severity failure;
	assert RAM(3866) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(3866))))  severity failure;
	assert RAM(3867) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(3867))))  severity failure;
	assert RAM(3868) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3868))))  severity failure;
	assert RAM(3869) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(3869))))  severity failure;
	assert RAM(3870) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3870))))  severity failure;
	assert RAM(3871) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(3871))))  severity failure;
	assert RAM(3872) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(3872))))  severity failure;
	assert RAM(3873) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(3873))))  severity failure;
	assert RAM(3874) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(3874))))  severity failure;
	assert RAM(3875) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(3875))))  severity failure;
	assert RAM(3876) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(3876))))  severity failure;
	assert RAM(3877) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(3877))))  severity failure;
	assert RAM(3878) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(3878))))  severity failure;
	assert RAM(3879) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(3879))))  severity failure;
	assert RAM(3880) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(3880))))  severity failure;
	assert RAM(3881) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(3881))))  severity failure;
	assert RAM(3882) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(3882))))  severity failure;
	assert RAM(3883) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(3883))))  severity failure;
	assert RAM(3884) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(3884))))  severity failure;
	assert RAM(3885) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(3885))))  severity failure;
	assert RAM(3886) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(3886))))  severity failure;
	assert RAM(3887) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(3887))))  severity failure;
	assert RAM(3888) = std_logic_vector(to_unsigned(220, 8)) report "TEST FALLITO (WORKING ZONE). Expected  220  found " & integer'image(to_integer(unsigned(RAM(3888))))  severity failure;
	assert RAM(3889) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(3889))))  severity failure;
	assert RAM(3890) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(3890))))  severity failure;
	assert RAM(3891) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(3891))))  severity failure;
	assert RAM(3892) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(3892))))  severity failure;
	assert RAM(3893) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(3893))))  severity failure;
	assert RAM(3894) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(3894))))  severity failure;
	assert RAM(3895) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(3895))))  severity failure;
	assert RAM(3896) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(3896))))  severity failure;
	assert RAM(3897) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(3897))))  severity failure;
	assert RAM(3898) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(3898))))  severity failure;
	assert RAM(3899) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(3899))))  severity failure;
	assert RAM(3900) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(3900))))  severity failure;
	assert RAM(3901) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(3901))))  severity failure;
	assert RAM(3902) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(3902))))  severity failure;
	assert RAM(3903) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(3903))))  severity failure;
	assert RAM(3904) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(3904))))  severity failure;
	assert RAM(3905) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(3905))))  severity failure;
	assert RAM(3906) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(3906))))  severity failure;
	assert RAM(3907) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(3907))))  severity failure;
	assert RAM(3908) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(3908))))  severity failure;
	assert RAM(3909) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(3909))))  severity failure;
	assert RAM(3910) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(3910))))  severity failure;
	assert RAM(3911) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(3911))))  severity failure;
	assert RAM(3912) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(3912))))  severity failure;
	assert RAM(3913) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(3913))))  severity failure;
	assert RAM(3914) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(3914))))  severity failure;
	assert RAM(3915) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(3915))))  severity failure;
	assert RAM(3916) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(3916))))  severity failure;
	assert RAM(3917) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(3917))))  severity failure;
	assert RAM(3918) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(3918))))  severity failure;
	assert RAM(3919) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(3919))))  severity failure;
	assert RAM(3920) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(3920))))  severity failure;
	assert RAM(3921) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(3921))))  severity failure;
	assert RAM(3922) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(3922))))  severity failure;
	assert RAM(3923) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(3923))))  severity failure;
	assert RAM(3924) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(3924))))  severity failure;
	assert RAM(3925) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(3925))))  severity failure;
	assert RAM(3926) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(3926))))  severity failure;
	assert RAM(3927) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(3927))))  severity failure;
	assert RAM(3928) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(3928))))  severity failure;
	assert RAM(3929) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(3929))))  severity failure;
	assert RAM(3930) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(3930))))  severity failure;
	assert RAM(3931) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(3931))))  severity failure;
	assert RAM(3932) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(3932))))  severity failure;
	assert RAM(3933) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(3933))))  severity failure;
	assert RAM(3934) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(3934))))  severity failure;
	assert RAM(3935) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(3935))))  severity failure;
	assert RAM(3936) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(3936))))  severity failure;
	assert RAM(3937) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(3937))))  severity failure;
	assert RAM(3938) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(3938))))  severity failure;
	assert RAM(3939) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(3939))))  severity failure;
	assert RAM(3940) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(3940))))  severity failure;
	assert RAM(3941) = std_logic_vector(to_unsigned(224, 8)) report "TEST FALLITO (WORKING ZONE). Expected  224  found " & integer'image(to_integer(unsigned(RAM(3941))))  severity failure;
	assert RAM(3942) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(3942))))  severity failure;
	assert RAM(3943) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(3943))))  severity failure;
	assert RAM(3944) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(3944))))  severity failure;
	assert RAM(3945) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3945))))  severity failure;
	assert RAM(3946) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(3946))))  severity failure;
	assert RAM(3947) = std_logic_vector(to_unsigned(41, 8)) report "TEST FALLITO (WORKING ZONE). Expected  41  found " & integer'image(to_integer(unsigned(RAM(3947))))  severity failure;
	assert RAM(3948) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(3948))))  severity failure;
	assert RAM(3949) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(3949))))  severity failure;
	assert RAM(3950) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(3950))))  severity failure;
	assert RAM(3951) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(3951))))  severity failure;
	assert RAM(3952) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(3952))))  severity failure;
	assert RAM(3953) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(3953))))  severity failure;
	assert RAM(3954) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(3954))))  severity failure;
	assert RAM(3955) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(3955))))  severity failure;
	assert RAM(3956) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(3956))))  severity failure;
	assert RAM(3957) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(3957))))  severity failure;
	assert RAM(3958) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(3958))))  severity failure;
	assert RAM(3959) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(3959))))  severity failure;
	assert RAM(3960) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(3960))))  severity failure;
	assert RAM(3961) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(3961))))  severity failure;
	assert RAM(3962) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(3962))))  severity failure;
	assert RAM(3963) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(3963))))  severity failure;
	assert RAM(3964) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(3964))))  severity failure;
	assert RAM(3965) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(3965))))  severity failure;
	assert RAM(3966) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(3966))))  severity failure;
	assert RAM(3967) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(3967))))  severity failure;
	assert RAM(3968) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(3968))))  severity failure;
	assert RAM(3969) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(3969))))  severity failure;
	assert RAM(3970) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(3970))))  severity failure;
	assert RAM(3971) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(3971))))  severity failure;
	assert RAM(3972) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(3972))))  severity failure;
	assert RAM(3973) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(3973))))  severity failure;
	assert RAM(3974) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(3974))))  severity failure;
	assert RAM(3975) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(3975))))  severity failure;
	assert RAM(3976) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(3976))))  severity failure;
	assert RAM(3977) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(3977))))  severity failure;
	assert RAM(3978) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3978))))  severity failure;
	assert RAM(3979) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(3979))))  severity failure;
	assert RAM(3980) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(3980))))  severity failure;
	assert RAM(3981) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(3981))))  severity failure;
	assert RAM(3982) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(3982))))  severity failure;
	assert RAM(3983) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(3983))))  severity failure;
	assert RAM(3984) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(3984))))  severity failure;
	assert RAM(3985) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(3985))))  severity failure;
	assert RAM(3986) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(3986))))  severity failure;
	assert RAM(3987) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(3987))))  severity failure;
	assert RAM(3988) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(3988))))  severity failure;
	assert RAM(3989) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(3989))))  severity failure;
	assert RAM(3990) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(3990))))  severity failure;
	assert RAM(3991) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(3991))))  severity failure;
	assert RAM(3992) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(3992))))  severity failure;
	assert RAM(3993) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(3993))))  severity failure;
	assert RAM(3994) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(3994))))  severity failure;
	assert RAM(3995) = std_logic_vector(to_unsigned(144, 8)) report "TEST FALLITO (WORKING ZONE). Expected  144  found " & integer'image(to_integer(unsigned(RAM(3995))))  severity failure;
	assert RAM(3996) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(3996))))  severity failure;
	assert RAM(3997) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(3997))))  severity failure;
	assert RAM(3998) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(3998))))  severity failure;
	assert RAM(3999) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(3999))))  severity failure;
	assert RAM(4000) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(4000))))  severity failure;
	assert RAM(4001) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(4001))))  severity failure;
	assert RAM(4002) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(4002))))  severity failure;
	assert RAM(4003) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(4003))))  severity failure;
	assert RAM(4004) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(4004))))  severity failure;
	assert RAM(4005) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(4005))))  severity failure;
	assert RAM(4006) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(4006))))  severity failure;
	assert RAM(4007) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(4007))))  severity failure;
	assert RAM(4008) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(4008))))  severity failure;
	assert RAM(4009) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(4009))))  severity failure;
	assert RAM(4010) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(4010))))  severity failure;
	assert RAM(4011) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(4011))))  severity failure;
	assert RAM(4012) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(4012))))  severity failure;
	assert RAM(4013) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(4013))))  severity failure;
	assert RAM(4014) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(4014))))  severity failure;
	assert RAM(4015) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(4015))))  severity failure;
	assert RAM(4016) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(4016))))  severity failure;
	assert RAM(4017) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(4017))))  severity failure;
	assert RAM(4018) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(4018))))  severity failure;
	assert RAM(4019) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(4019))))  severity failure;
	assert RAM(4020) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(4020))))  severity failure;
	assert RAM(4021) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(4021))))  severity failure;
	assert RAM(4022) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(4022))))  severity failure;
	assert RAM(4023) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(4023))))  severity failure;
	assert RAM(4024) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(4024))))  severity failure;
	assert RAM(4025) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(4025))))  severity failure;
	assert RAM(4026) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(4026))))  severity failure;
	assert RAM(4027) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(4027))))  severity failure;
	assert RAM(4028) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(4028))))  severity failure;
	assert RAM(4029) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(4029))))  severity failure;
	assert RAM(4030) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(4030))))  severity failure;
	assert RAM(4031) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(4031))))  severity failure;
	assert RAM(4032) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(4032))))  severity failure;
	assert RAM(4033) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(4033))))  severity failure;
	assert RAM(4034) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(4034))))  severity failure;
	assert RAM(4035) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(4035))))  severity failure;
	assert RAM(4036) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(4036))))  severity failure;
	assert RAM(4037) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(4037))))  severity failure;
	assert RAM(4038) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(4038))))  severity failure;
	assert RAM(4039) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(4039))))  severity failure;
	assert RAM(4040) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(4040))))  severity failure;
	assert RAM(4041) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(4041))))  severity failure;
	assert RAM(4042) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(4042))))  severity failure;
	assert RAM(4043) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(4043))))  severity failure;
	assert RAM(4044) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(4044))))  severity failure;
	assert RAM(4045) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(4045))))  severity failure;
	assert RAM(4046) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(4046))))  severity failure;
	assert RAM(4047) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(4047))))  severity failure;
	assert RAM(4048) = std_logic_vector(to_unsigned(60, 8)) report "TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM(4048))))  severity failure;
	assert RAM(4049) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(4049))))  severity failure;
	assert RAM(4050) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(4050))))  severity failure;
	assert RAM(4051) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(4051))))  severity failure;
	assert RAM(4052) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(4052))))  severity failure;
	assert RAM(4053) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(4053))))  severity failure;
	assert RAM(4054) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(4054))))  severity failure;
	assert RAM(4055) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(4055))))  severity failure;
	assert RAM(4056) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(4056))))  severity failure;
	assert RAM(4057) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(4057))))  severity failure;
	assert RAM(4058) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(4058))))  severity failure;
	assert RAM(4059) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(4059))))  severity failure;
	assert RAM(4060) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(4060))))  severity failure;
	assert RAM(4061) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(4061))))  severity failure;
	assert RAM(4062) = std_logic_vector(to_unsigned(59, 8)) report "TEST FALLITO (WORKING ZONE). Expected  59  found " & integer'image(to_integer(unsigned(RAM(4062))))  severity failure;
	assert RAM(4063) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(4063))))  severity failure;
	assert RAM(4064) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(4064))))  severity failure;
	assert RAM(4065) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(4065))))  severity failure;
	assert RAM(4066) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(4066))))  severity failure;
	assert RAM(4067) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(4067))))  severity failure;
	assert RAM(4068) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(4068))))  severity failure;
	assert RAM(4069) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(4069))))  severity failure;
	assert RAM(4070) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(4070))))  severity failure;
	assert RAM(4071) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(4071))))  severity failure;
	assert RAM(4072) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(4072))))  severity failure;
	assert RAM(4073) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(4073))))  severity failure;
	assert RAM(4074) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(4074))))  severity failure;
	assert RAM(4075) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(4075))))  severity failure;
	assert RAM(4076) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(4076))))  severity failure;
	assert RAM(4077) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(4077))))  severity failure;
	assert RAM(4078) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(4078))))  severity failure;
	assert RAM(4079) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(4079))))  severity failure;
	assert RAM(4080) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(4080))))  severity failure;
	assert RAM(4081) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(4081))))  severity failure;
	assert RAM(4082) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(4082))))  severity failure;
	assert RAM(4083) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(4083))))  severity failure;
	assert RAM(4084) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(4084))))  severity failure;
	assert RAM(4085) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(4085))))  severity failure;
	assert RAM(4086) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(4086))))  severity failure;
	assert RAM(4087) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(4087))))  severity failure;
	assert RAM(4088) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(4088))))  severity failure;
	assert RAM(4089) = std_logic_vector(to_unsigned(121, 8)) report "TEST FALLITO (WORKING ZONE). Expected  121  found " & integer'image(to_integer(unsigned(RAM(4089))))  severity failure;
	assert RAM(4090) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(4090))))  severity failure;
	assert RAM(4091) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(4091))))  severity failure;
	assert RAM(4092) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(4092))))  severity failure;
	assert RAM(4093) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(4093))))  severity failure;
	assert RAM(4094) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(4094))))  severity failure;
	assert RAM(4095) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(4095))))  severity failure;
	assert RAM(4096) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(4096))))  severity failure;
	assert RAM(4097) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(4097))))  severity failure;
	assert RAM(4098) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(4098))))  severity failure;
	assert RAM(4099) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(4099))))  severity failure;
	assert RAM(4100) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(4100))))  severity failure;
	assert RAM(4101) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(4101))))  severity failure;
	assert RAM(4102) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(4102))))  severity failure;
	assert RAM(4103) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(4103))))  severity failure;
	assert RAM(4104) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(4104))))  severity failure;
	assert RAM(4105) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(4105))))  severity failure;
	assert RAM(4106) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(4106))))  severity failure;
	assert RAM(4107) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(4107))))  severity failure;
	assert RAM(4108) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(4108))))  severity failure;
	assert RAM(4109) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(4109))))  severity failure;
	assert RAM(4110) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(4110))))  severity failure;
	assert RAM(4111) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(4111))))  severity failure;
	assert RAM(4112) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(4112))))  severity failure;
	assert RAM(4113) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(4113))))  severity failure;
	assert RAM(4114) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(4114))))  severity failure;
	assert RAM(4115) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(4115))))  severity failure;
	assert RAM(4116) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(4116))))  severity failure;
	assert RAM(4117) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(4117))))  severity failure;
	assert RAM(4118) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(4118))))  severity failure;
	assert RAM(4119) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(4119))))  severity failure;
	assert RAM(4120) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(4120))))  severity failure;
	assert RAM(4121) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(4121))))  severity failure;
	assert RAM(4122) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(4122))))  severity failure;
	assert RAM(4123) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(4123))))  severity failure;
	assert RAM(4124) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(4124))))  severity failure;
	assert RAM(4125) = std_logic_vector(to_unsigned(162, 8)) report "TEST FALLITO (WORKING ZONE). Expected  162  found " & integer'image(to_integer(unsigned(RAM(4125))))  severity failure;
	assert RAM(4126) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(4126))))  severity failure;
	assert RAM(4127) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(4127))))  severity failure;
	assert RAM(4128) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(4128))))  severity failure;
	assert RAM(4129) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(4129))))  severity failure;
	assert RAM(4130) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(4130))))  severity failure;
	assert RAM(4131) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(4131))))  severity failure;
	assert RAM(4132) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(4132))))  severity failure;
	assert RAM(4133) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(4133))))  severity failure;
	assert RAM(4134) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(4134))))  severity failure;
	assert RAM(4135) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(4135))))  severity failure;
	assert RAM(4136) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(4136))))  severity failure;
	assert RAM(4137) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(4137))))  severity failure;
	assert RAM(4138) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(4138))))  severity failure;
	assert RAM(4139) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(4139))))  severity failure;
	assert RAM(4140) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(4140))))  severity failure;
	assert RAM(4141) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(4141))))  severity failure;
	assert RAM(4142) = std_logic_vector(to_unsigned(110, 8)) report "TEST FALLITO (WORKING ZONE). Expected  110  found " & integer'image(to_integer(unsigned(RAM(4142))))  severity failure;
	assert RAM(4143) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(4143))))  severity failure;
	assert RAM(4144) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(4144))))  severity failure;
	assert RAM(4145) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(4145))))  severity failure;
	assert RAM(4146) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(4146))))  severity failure;
	assert RAM(4147) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(4147))))  severity failure;
	assert RAM(4148) = std_logic_vector(to_unsigned(127, 8)) report "TEST FALLITO (WORKING ZONE). Expected  127  found " & integer'image(to_integer(unsigned(RAM(4148))))  severity failure;
	assert RAM(4149) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(4149))))  severity failure;
	assert RAM(4150) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(4150))))  severity failure;
	assert RAM(4151) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(4151))))  severity failure;
	assert RAM(4152) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(4152))))  severity failure;
	assert RAM(4153) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(4153))))  severity failure;
	assert RAM(4154) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(4154))))  severity failure;
	assert RAM(4155) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(4155))))  severity failure;
	assert RAM(4156) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(4156))))  severity failure;
	assert RAM(4157) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(4157))))  severity failure;
	assert RAM(4158) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(4158))))  severity failure;
	assert RAM(4159) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(4159))))  severity failure;
	assert RAM(4160) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(4160))))  severity failure;
	assert RAM(4161) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(4161))))  severity failure;
	assert RAM(4162) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(4162))))  severity failure;
	assert RAM(4163) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(4163))))  severity failure;
	assert RAM(4164) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(4164))))  severity failure;
	assert RAM(4165) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(4165))))  severity failure;
	assert RAM(4166) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(4166))))  severity failure;
	assert RAM(4167) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(4167))))  severity failure;
	assert RAM(4168) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(4168))))  severity failure;
	assert RAM(4169) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(4169))))  severity failure;
	assert RAM(4170) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(4170))))  severity failure;
	assert RAM(4171) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(4171))))  severity failure;
	assert RAM(4172) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(4172))))  severity failure;
	assert RAM(4173) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(4173))))  severity failure;
	assert RAM(4174) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(4174))))  severity failure;
	assert RAM(4175) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(4175))))  severity failure;
	assert RAM(4176) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(4176))))  severity failure;
	assert RAM(4177) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(4177))))  severity failure;
	assert RAM(4178) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(4178))))  severity failure;
	assert RAM(4179) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(4179))))  severity failure;
	assert RAM(4180) = std_logic_vector(to_unsigned(194, 8)) report "TEST FALLITO (WORKING ZONE). Expected  194  found " & integer'image(to_integer(unsigned(RAM(4180))))  severity failure;
	assert RAM(4181) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(4181))))  severity failure;
	assert RAM(4182) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(4182))))  severity failure;
	assert RAM(4183) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(4183))))  severity failure;
	assert RAM(4184) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(4184))))  severity failure;
	assert RAM(4185) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(4185))))  severity failure;
	assert RAM(4186) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(4186))))  severity failure;
	assert RAM(4187) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(4187))))  severity failure;
	assert RAM(4188) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(4188))))  severity failure;
	assert RAM(4189) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(4189))))  severity failure;
	assert RAM(4190) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(4190))))  severity failure;
	assert RAM(4191) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(4191))))  severity failure;
	assert RAM(4192) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(4192))))  severity failure;
	assert RAM(4193) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(4193))))  severity failure;
	assert RAM(4194) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(4194))))  severity failure;
	assert RAM(4195) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(4195))))  severity failure;
	assert RAM(4196) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(4196))))  severity failure;
	assert RAM(4197) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(4197))))  severity failure;
	assert RAM(4198) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(4198))))  severity failure;
	assert RAM(4199) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(4199))))  severity failure;
	assert RAM(4200) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(4200))))  severity failure;
	assert RAM(4201) = std_logic_vector(to_unsigned(89, 8)) report "TEST FALLITO (WORKING ZONE). Expected  89  found " & integer'image(to_integer(unsigned(RAM(4201))))  severity failure;
	assert RAM(4202) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(4202))))  severity failure;
	assert RAM(4203) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(4203))))  severity failure;
	assert RAM(4204) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(4204))))  severity failure;
	assert RAM(4205) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(4205))))  severity failure;
	assert RAM(4206) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(4206))))  severity failure;
	assert RAM(4207) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(4207))))  severity failure;
	assert RAM(4208) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(4208))))  severity failure;
	assert RAM(4209) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(4209))))  severity failure;
	assert RAM(4210) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(4210))))  severity failure;
	assert RAM(4211) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(4211))))  severity failure;
	assert RAM(4212) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(4212))))  severity failure;
	assert RAM(4213) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(4213))))  severity failure;
	assert RAM(4214) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(4214))))  severity failure;
	assert RAM(4215) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(4215))))  severity failure;
	assert RAM(4216) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(4216))))  severity failure;
	assert RAM(4217) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(4217))))  severity failure;
	assert RAM(4218) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(4218))))  severity failure;
	assert RAM(4219) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(4219))))  severity failure;
	assert RAM(4220) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(4220))))  severity failure;
	assert RAM(4221) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(4221))))  severity failure;
	assert RAM(4222) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(4222))))  severity failure;
	assert RAM(4223) = std_logic_vector(to_unsigned(168, 8)) report "TEST FALLITO (WORKING ZONE). Expected  168  found " & integer'image(to_integer(unsigned(RAM(4223))))  severity failure;
	assert RAM(4224) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(4224))))  severity failure;
	assert RAM(4225) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(4225))))  severity failure;
	assert RAM(4226) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(4226))))  severity failure;
	assert RAM(4227) = std_logic_vector(to_unsigned(75, 8)) report "TEST FALLITO (WORKING ZONE). Expected  75  found " & integer'image(to_integer(unsigned(RAM(4227))))  severity failure;
	assert RAM(4228) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(4228))))  severity failure;
	assert RAM(4229) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(4229))))  severity failure;
	assert RAM(4230) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(4230))))  severity failure;
	assert RAM(4231) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(4231))))  severity failure;
	assert RAM(4232) = std_logic_vector(to_unsigned(49, 8)) report "TEST FALLITO (WORKING ZONE). Expected  49  found " & integer'image(to_integer(unsigned(RAM(4232))))  severity failure;
	assert RAM(4233) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(4233))))  severity failure;
	assert RAM(4234) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(4234))))  severity failure;
	assert RAM(4235) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(4235))))  severity failure;
	assert RAM(4236) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(4236))))  severity failure;
	assert RAM(4237) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(4237))))  severity failure;
	assert RAM(4238) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(4238))))  severity failure;
	assert RAM(4239) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(4239))))  severity failure;
	assert RAM(4240) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(4240))))  severity failure;
	assert RAM(4241) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(4241))))  severity failure;
	assert RAM(4242) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(4242))))  severity failure;
	assert RAM(4243) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(4243))))  severity failure;
	assert RAM(4244) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(4244))))  severity failure;
	assert RAM(4245) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(4245))))  severity failure;
	assert RAM(4246) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(4246))))  severity failure;
	assert RAM(4247) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(4247))))  severity failure;
	assert RAM(4248) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(4248))))  severity failure;
	assert RAM(4249) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(4249))))  severity failure;
	assert RAM(4250) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(4250))))  severity failure;
	assert RAM(4251) = std_logic_vector(to_unsigned(138, 8)) report "TEST FALLITO (WORKING ZONE). Expected  138  found " & integer'image(to_integer(unsigned(RAM(4251))))  severity failure;
	assert RAM(4252) = std_logic_vector(to_unsigned(204, 8)) report "TEST FALLITO (WORKING ZONE). Expected  204  found " & integer'image(to_integer(unsigned(RAM(4252))))  severity failure;
	assert RAM(4253) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(4253))))  severity failure;
	assert RAM(4254) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(4254))))  severity failure;
	assert RAM(4255) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(4255))))  severity failure;
	assert RAM(4256) = std_logic_vector(to_unsigned(57, 8)) report "TEST FALLITO (WORKING ZONE). Expected  57  found " & integer'image(to_integer(unsigned(RAM(4256))))  severity failure;
	assert RAM(4257) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(4257))))  severity failure;
	assert RAM(4258) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(4258))))  severity failure;
	assert RAM(4259) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(4259))))  severity failure;
	assert RAM(4260) = std_logic_vector(to_unsigned(125, 8)) report "TEST FALLITO (WORKING ZONE). Expected  125  found " & integer'image(to_integer(unsigned(RAM(4260))))  severity failure;
	assert RAM(4261) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(4261))))  severity failure;
	assert RAM(4262) = std_logic_vector(to_unsigned(16, 8)) report "TEST FALLITO (WORKING ZONE). Expected  16  found " & integer'image(to_integer(unsigned(RAM(4262))))  severity failure;
	assert RAM(4263) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(4263))))  severity failure;
	assert RAM(4264) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(4264))))  severity failure;
	assert RAM(4265) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(4265))))  severity failure;
	assert RAM(4266) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(4266))))  severity failure;
	assert RAM(4267) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(4267))))  severity failure;
	assert RAM(4268) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(4268))))  severity failure;
	assert RAM(4269) = std_logic_vector(to_unsigned(39, 8)) report "TEST FALLITO (WORKING ZONE). Expected  39  found " & integer'image(to_integer(unsigned(RAM(4269))))  severity failure;
	assert RAM(4270) = std_logic_vector(to_unsigned(218, 8)) report "TEST FALLITO (WORKING ZONE). Expected  218  found " & integer'image(to_integer(unsigned(RAM(4270))))  severity failure;
	assert RAM(4271) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(4271))))  severity failure;
	assert RAM(4272) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(4272))))  severity failure;
	assert RAM(4273) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(4273))))  severity failure;
	assert RAM(4274) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(4274))))  severity failure;
	assert RAM(4275) = std_logic_vector(to_unsigned(183, 8)) report "TEST FALLITO (WORKING ZONE). Expected  183  found " & integer'image(to_integer(unsigned(RAM(4275))))  severity failure;
	assert RAM(4276) = std_logic_vector(to_unsigned(195, 8)) report "TEST FALLITO (WORKING ZONE). Expected  195  found " & integer'image(to_integer(unsigned(RAM(4276))))  severity failure;
	assert RAM(4277) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(4277))))  severity failure;
	assert RAM(4278) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(4278))))  severity failure;
	assert RAM(4279) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(4279))))  severity failure;
	assert RAM(4280) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(4280))))  severity failure;
	assert RAM(4281) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(4281))))  severity failure;
	assert RAM(4282) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(4282))))  severity failure;
	assert RAM(4283) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(4283))))  severity failure;
	assert RAM(4284) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(4284))))  severity failure;
	assert RAM(4285) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(4285))))  severity failure;
	assert RAM(4286) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(4286))))  severity failure;
	assert RAM(4287) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(4287))))  severity failure;
	assert RAM(4288) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(4288))))  severity failure;
	assert RAM(4289) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(4289))))  severity failure;
	assert RAM(4290) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(4290))))  severity failure;
	assert RAM(4291) = std_logic_vector(to_unsigned(145, 8)) report "TEST FALLITO (WORKING ZONE). Expected  145  found " & integer'image(to_integer(unsigned(RAM(4291))))  severity failure;
	assert RAM(4292) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(4292))))  severity failure;
	assert RAM(4293) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(4293))))  severity failure;
	assert RAM(4294) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(4294))))  severity failure;
	assert RAM(4295) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(4295))))  severity failure;
	assert RAM(4296) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(4296))))  severity failure;
	assert RAM(4297) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(4297))))  severity failure;
	assert RAM(4298) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(4298))))  severity failure;
	assert RAM(4299) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(4299))))  severity failure;
	assert RAM(4300) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(4300))))  severity failure;
	assert RAM(4301) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(4301))))  severity failure;
	assert RAM(4302) = std_logic_vector(to_unsigned(134, 8)) report "TEST FALLITO (WORKING ZONE). Expected  134  found " & integer'image(to_integer(unsigned(RAM(4302))))  severity failure;
	assert RAM(4303) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(4303))))  severity failure;
	assert RAM(4304) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(4304))))  severity failure;
	assert RAM(4305) = std_logic_vector(to_unsigned(129, 8)) report "TEST FALLITO (WORKING ZONE). Expected  129  found " & integer'image(to_integer(unsigned(RAM(4305))))  severity failure;
	assert RAM(4306) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(4306))))  severity failure;
	assert RAM(4307) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(4307))))  severity failure;
	assert RAM(4308) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(4308))))  severity failure;
	assert RAM(4309) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(4309))))  severity failure;
	assert RAM(4310) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(4310))))  severity failure;
	assert RAM(4311) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(4311))))  severity failure;
	assert RAM(4312) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(4312))))  severity failure;
	assert RAM(4313) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(4313))))  severity failure;
	assert RAM(4314) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(4314))))  severity failure;
	assert RAM(4315) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(4315))))  severity failure;
	assert RAM(4316) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(4316))))  severity failure;
	assert RAM(4317) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(4317))))  severity failure;
	assert RAM(4318) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(4318))))  severity failure;
	assert RAM(4319) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(4319))))  severity failure;
	assert RAM(4320) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(4320))))  severity failure;
	assert RAM(4321) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(4321))))  severity failure;
	assert RAM(4322) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(4322))))  severity failure;
	assert RAM(4323) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(4323))))  severity failure;
	assert RAM(4324) = std_logic_vector(to_unsigned(199, 8)) report "TEST FALLITO (WORKING ZONE). Expected  199  found " & integer'image(to_integer(unsigned(RAM(4324))))  severity failure;
	assert RAM(4325) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(4325))))  severity failure;
	assert RAM(4326) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(4326))))  severity failure;
	assert RAM(4327) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(4327))))  severity failure;
	assert RAM(4328) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(4328))))  severity failure;
	assert RAM(4329) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(4329))))  severity failure;
	assert RAM(4330) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(4330))))  severity failure;
	assert RAM(4331) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(4331))))  severity failure;
	assert RAM(4332) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(4332))))  severity failure;
	assert RAM(4333) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(4333))))  severity failure;
	assert RAM(4334) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(4334))))  severity failure;
	assert RAM(4335) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(4335))))  severity failure;
	assert RAM(4336) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(4336))))  severity failure;
	assert RAM(4337) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(4337))))  severity failure;
	assert RAM(4338) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(4338))))  severity failure;
	assert RAM(4339) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(4339))))  severity failure;
	assert RAM(4340) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(4340))))  severity failure;
	assert RAM(4341) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(4341))))  severity failure;
	assert RAM(4342) = std_logic_vector(to_unsigned(87, 8)) report "TEST FALLITO (WORKING ZONE). Expected  87  found " & integer'image(to_integer(unsigned(RAM(4342))))  severity failure;
	assert RAM(4343) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(4343))))  severity failure;
	assert RAM(4344) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(4344))))  severity failure;
	assert RAM(4345) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(4345))))  severity failure;
	assert RAM(4346) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(4346))))  severity failure;
	assert RAM(4347) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(4347))))  severity failure;
	assert RAM(4348) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(4348))))  severity failure;
	assert RAM(4349) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(4349))))  severity failure;
	assert RAM(4350) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(4350))))  severity failure;
	assert RAM(4351) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(4351))))  severity failure;
	assert RAM(4352) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(4352))))  severity failure;
	assert RAM(4353) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(4353))))  severity failure;
	assert RAM(4354) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(4354))))  severity failure;
	assert RAM(4355) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(4355))))  severity failure;
	assert RAM(4356) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(4356))))  severity failure;
	assert RAM(4357) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(4357))))  severity failure;
	assert RAM(4358) = std_logic_vector(to_unsigned(241, 8)) report "TEST FALLITO (WORKING ZONE). Expected  241  found " & integer'image(to_integer(unsigned(RAM(4358))))  severity failure;
	assert RAM(4359) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(4359))))  severity failure;
	assert RAM(4360) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(4360))))  severity failure;
	assert RAM(4361) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(4361))))  severity failure;
	assert RAM(4362) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(4362))))  severity failure;
	assert RAM(4363) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(4363))))  severity failure;
	assert RAM(4364) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(4364))))  severity failure;
	assert RAM(4365) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(4365))))  severity failure;
	assert RAM(4366) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(4366))))  severity failure;
	assert RAM(4367) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(4367))))  severity failure;
	assert RAM(4368) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(4368))))  severity failure;
	assert RAM(4369) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(4369))))  severity failure;
	assert RAM(4370) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(4370))))  severity failure;
	assert RAM(4371) = std_logic_vector(to_unsigned(143, 8)) report "TEST FALLITO (WORKING ZONE). Expected  143  found " & integer'image(to_integer(unsigned(RAM(4371))))  severity failure;
	assert RAM(4372) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(4372))))  severity failure;
	assert RAM(4373) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(4373))))  severity failure;
	assert RAM(4374) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(4374))))  severity failure;
	assert RAM(4375) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(4375))))  severity failure;
	assert RAM(4376) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(4376))))  severity failure;
	assert RAM(4377) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(4377))))  severity failure;
	assert RAM(4378) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(4378))))  severity failure;
	assert RAM(4379) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(4379))))  severity failure;
	assert RAM(4380) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(4380))))  severity failure;
	assert RAM(4381) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(4381))))  severity failure;
	assert RAM(4382) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(4382))))  severity failure;
	assert RAM(4383) = std_logic_vector(to_unsigned(31, 8)) report "TEST FALLITO (WORKING ZONE). Expected  31  found " & integer'image(to_integer(unsigned(RAM(4383))))  severity failure;
	assert RAM(4384) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(4384))))  severity failure;
	assert RAM(4385) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(4385))))  severity failure;
	assert RAM(4386) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(4386))))  severity failure;
	assert RAM(4387) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(4387))))  severity failure;
	assert RAM(4388) = std_logic_vector(to_unsigned(119, 8)) report "TEST FALLITO (WORKING ZONE). Expected  119  found " & integer'image(to_integer(unsigned(RAM(4388))))  severity failure;
	assert RAM(4389) = std_logic_vector(to_unsigned(171, 8)) report "TEST FALLITO (WORKING ZONE). Expected  171  found " & integer'image(to_integer(unsigned(RAM(4389))))  severity failure;
	assert RAM(4390) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(4390))))  severity failure;
	assert RAM(4391) = std_logic_vector(to_unsigned(78, 8)) report "TEST FALLITO (WORKING ZONE). Expected  78  found " & integer'image(to_integer(unsigned(RAM(4391))))  severity failure;
	assert RAM(4392) = std_logic_vector(to_unsigned(13, 8)) report "TEST FALLITO (WORKING ZONE). Expected  13  found " & integer'image(to_integer(unsigned(RAM(4392))))  severity failure;
	assert RAM(4393) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(4393))))  severity failure;
	assert RAM(4394) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(4394))))  severity failure;
	assert RAM(4395) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(4395))))  severity failure;
	assert RAM(4396) = std_logic_vector(to_unsigned(104, 8)) report "TEST FALLITO (WORKING ZONE). Expected  104  found " & integer'image(to_integer(unsigned(RAM(4396))))  severity failure;
	assert RAM(4397) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(4397))))  severity failure;
	assert RAM(4398) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(4398))))  severity failure;
	assert RAM(4399) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(4399))))  severity failure;
	assert RAM(4400) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(4400))))  severity failure;
	assert RAM(4401) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(4401))))  severity failure;
	assert RAM(4402) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(4402))))  severity failure;
	assert RAM(4403) = std_logic_vector(to_unsigned(38, 8)) report "TEST FALLITO (WORKING ZONE). Expected  38  found " & integer'image(to_integer(unsigned(RAM(4403))))  severity failure;
	assert RAM(4404) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(4404))))  severity failure;
	assert RAM(4405) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(4405))))  severity failure;
	assert RAM(4406) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(4406))))  severity failure;
	assert RAM(4407) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(4407))))  severity failure;
	assert RAM(4408) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(4408))))  severity failure;
	assert RAM(4409) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(4409))))  severity failure;
	assert RAM(4410) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(4410))))  severity failure;
	assert RAM(4411) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(4411))))  severity failure;
	assert RAM(4412) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(4412))))  severity failure;
	assert RAM(4413) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(4413))))  severity failure;
	assert RAM(4414) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(4414))))  severity failure;
	assert RAM(4415) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(4415))))  severity failure;
	assert RAM(4416) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(4416))))  severity failure;
	assert RAM(4417) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(4417))))  severity failure;
	assert RAM(4418) = std_logic_vector(to_unsigned(187, 8)) report "TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM(4418))))  severity failure;
	assert RAM(4419) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(4419))))  severity failure;
	assert RAM(4420) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(4420))))  severity failure;
	assert RAM(4421) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(4421))))  severity failure;
	assert RAM(4422) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(4422))))  severity failure;
	assert RAM(4423) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(4423))))  severity failure;
	assert RAM(4424) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(4424))))  severity failure;
	assert RAM(4425) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(4425))))  severity failure;
	assert RAM(4426) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(4426))))  severity failure;
	assert RAM(4427) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(4427))))  severity failure;
	assert RAM(4428) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(4428))))  severity failure;
	assert RAM(4429) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(4429))))  severity failure;
	assert RAM(4430) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(4430))))  severity failure;
	assert RAM(4431) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(4431))))  severity failure;
	assert RAM(4432) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(4432))))  severity failure;
	assert RAM(4433) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(4433))))  severity failure;
	assert RAM(4434) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(4434))))  severity failure;
	assert RAM(4435) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(4435))))  severity failure;
	assert RAM(4436) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(4436))))  severity failure;
	assert RAM(4437) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(4437))))  severity failure;
	assert RAM(4438) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(4438))))  severity failure;
	assert RAM(4439) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(4439))))  severity failure;
	assert RAM(4440) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(4440))))  severity failure;
	assert RAM(4441) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(4441))))  severity failure;
	assert RAM(4442) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(4442))))  severity failure;
	assert RAM(4443) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(4443))))  severity failure;
	assert RAM(4444) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(4444))))  severity failure;
	assert RAM(4445) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(4445))))  severity failure;
	assert RAM(4446) = std_logic_vector(to_unsigned(253, 8)) report "TEST FALLITO (WORKING ZONE). Expected  253  found " & integer'image(to_integer(unsigned(RAM(4446))))  severity failure;
	assert RAM(4447) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(4447))))  severity failure;
	assert RAM(4448) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(4448))))  severity failure;
	assert RAM(4449) = std_logic_vector(to_unsigned(212, 8)) report "TEST FALLITO (WORKING ZONE). Expected  212  found " & integer'image(to_integer(unsigned(RAM(4449))))  severity failure;
	assert RAM(4450) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(4450))))  severity failure;
	assert RAM(4451) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(4451))))  severity failure;
	assert RAM(4452) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(4452))))  severity failure;
	assert RAM(4453) = std_logic_vector(to_unsigned(131, 8)) report "TEST FALLITO (WORKING ZONE). Expected  131  found " & integer'image(to_integer(unsigned(RAM(4453))))  severity failure;
	assert RAM(4454) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(4454))))  severity failure;
	assert RAM(4455) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(4455))))  severity failure;
	assert RAM(4456) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(4456))))  severity failure;
	assert RAM(4457) = std_logic_vector(to_unsigned(149, 8)) report "TEST FALLITO (WORKING ZONE). Expected  149  found " & integer'image(to_integer(unsigned(RAM(4457))))  severity failure;
	assert RAM(4458) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(4458))))  severity failure;
	assert RAM(4459) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(4459))))  severity failure;
	assert RAM(4460) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(4460))))  severity failure;
	assert RAM(4461) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(4461))))  severity failure;
	assert RAM(4462) = std_logic_vector(to_unsigned(85, 8)) report "TEST FALLITO (WORKING ZONE). Expected  85  found " & integer'image(to_integer(unsigned(RAM(4462))))  severity failure;
	assert RAM(4463) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(4463))))  severity failure;
	assert RAM(4464) = std_logic_vector(to_unsigned(150, 8)) report "TEST FALLITO (WORKING ZONE). Expected  150  found " & integer'image(to_integer(unsigned(RAM(4464))))  severity failure;
	assert RAM(4465) = std_logic_vector(to_unsigned(157, 8)) report "TEST FALLITO (WORKING ZONE). Expected  157  found " & integer'image(to_integer(unsigned(RAM(4465))))  severity failure;
	assert RAM(4466) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(4466))))  severity failure;
	assert RAM(4467) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(4467))))  severity failure;
	assert RAM(4468) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(4468))))  severity failure;
	assert RAM(4469) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(4469))))  severity failure;
	assert RAM(4470) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(4470))))  severity failure;
	assert RAM(4471) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(4471))))  severity failure;
	assert RAM(4472) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(4472))))  severity failure;
	assert RAM(4473) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(4473))))  severity failure;
	assert RAM(4474) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(4474))))  severity failure;
	assert RAM(4475) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(4475))))  severity failure;
	assert RAM(4476) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(4476))))  severity failure;
	assert RAM(4477) = std_logic_vector(to_unsigned(126, 8)) report "TEST FALLITO (WORKING ZONE). Expected  126  found " & integer'image(to_integer(unsigned(RAM(4477))))  severity failure;
	assert RAM(4478) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(4478))))  severity failure;
	assert RAM(4479) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(4479))))  severity failure;
	assert RAM(4480) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(4480))))  severity failure;
	assert RAM(4481) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(4481))))  severity failure;
	assert RAM(4482) = std_logic_vector(to_unsigned(37, 8)) report "TEST FALLITO (WORKING ZONE). Expected  37  found " & integer'image(to_integer(unsigned(RAM(4482))))  severity failure;
	assert RAM(4483) = std_logic_vector(to_unsigned(86, 8)) report "TEST FALLITO (WORKING ZONE). Expected  86  found " & integer'image(to_integer(unsigned(RAM(4483))))  severity failure;
	assert RAM(4484) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(4484))))  severity failure;
	assert RAM(4485) = std_logic_vector(to_unsigned(237, 8)) report "TEST FALLITO (WORKING ZONE). Expected  237  found " & integer'image(to_integer(unsigned(RAM(4485))))  severity failure;
	assert RAM(4486) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(4486))))  severity failure;
	assert RAM(4487) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(4487))))  severity failure;
	assert RAM(4488) = std_logic_vector(to_unsigned(35, 8)) report "TEST FALLITO (WORKING ZONE). Expected  35  found " & integer'image(to_integer(unsigned(RAM(4488))))  severity failure;
	assert RAM(4489) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(4489))))  severity failure;
	assert RAM(4490) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(4490))))  severity failure;
	assert RAM(4491) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(4491))))  severity failure;
	assert RAM(4492) = std_logic_vector(to_unsigned(73, 8)) report "TEST FALLITO (WORKING ZONE). Expected  73  found " & integer'image(to_integer(unsigned(RAM(4492))))  severity failure;
	assert RAM(4493) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(4493))))  severity failure;
	assert RAM(4494) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(4494))))  severity failure;
	assert RAM(4495) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(4495))))  severity failure;
	assert RAM(4496) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(4496))))  severity failure;
	assert RAM(4497) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(4497))))  severity failure;
	assert RAM(4498) = std_logic_vector(to_unsigned(249, 8)) report "TEST FALLITO (WORKING ZONE). Expected  249  found " & integer'image(to_integer(unsigned(RAM(4498))))  severity failure;
	assert RAM(4499) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(4499))))  severity failure;
	assert RAM(4500) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(4500))))  severity failure;
	assert RAM(4501) = std_logic_vector(to_unsigned(207, 8)) report "TEST FALLITO (WORKING ZONE). Expected  207  found " & integer'image(to_integer(unsigned(RAM(4501))))  severity failure;
	assert RAM(4502) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(4502))))  severity failure;
	assert RAM(4503) = std_logic_vector(to_unsigned(29, 8)) report "TEST FALLITO (WORKING ZONE). Expected  29  found " & integer'image(to_integer(unsigned(RAM(4503))))  severity failure;
	assert RAM(4504) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(4504))))  severity failure;
	assert RAM(4505) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(4505))))  severity failure;
	assert RAM(4506) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(4506))))  severity failure;
	assert RAM(4507) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(4507))))  severity failure;
	assert RAM(4508) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(4508))))  severity failure;
	assert RAM(4509) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(4509))))  severity failure;
	assert RAM(4510) = std_logic_vector(to_unsigned(99, 8)) report "TEST FALLITO (WORKING ZONE). Expected  99  found " & integer'image(to_integer(unsigned(RAM(4510))))  severity failure;
	assert RAM(4511) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(4511))))  severity failure;
	assert RAM(4512) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(4512))))  severity failure;
	assert RAM(4513) = std_logic_vector(to_unsigned(17, 8)) report "TEST FALLITO (WORKING ZONE). Expected  17  found " & integer'image(to_integer(unsigned(RAM(4513))))  severity failure;
	assert RAM(4514) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(4514))))  severity failure;
	assert RAM(4515) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(4515))))  severity failure;
	assert RAM(4516) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(4516))))  severity failure;
	assert RAM(4517) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(4517))))  severity failure;
	assert RAM(4518) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(4518))))  severity failure;
	assert RAM(4519) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(4519))))  severity failure;
	assert RAM(4520) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(4520))))  severity failure;
	assert RAM(4521) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(4521))))  severity failure;
	assert RAM(4522) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(4522))))  severity failure;
	assert RAM(4523) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(4523))))  severity failure;
	assert RAM(4524) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(4524))))  severity failure;
	assert RAM(4525) = std_logic_vector(to_unsigned(235, 8)) report "TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM(4525))))  severity failure;
	assert RAM(4526) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(4526))))  severity failure;
	assert RAM(4527) = std_logic_vector(to_unsigned(151, 8)) report "TEST FALLITO (WORKING ZONE). Expected  151  found " & integer'image(to_integer(unsigned(RAM(4527))))  severity failure;
	assert RAM(4528) = std_logic_vector(to_unsigned(69, 8)) report "TEST FALLITO (WORKING ZONE). Expected  69  found " & integer'image(to_integer(unsigned(RAM(4528))))  severity failure;
	assert RAM(4529) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(4529))))  severity failure;
	assert RAM(4530) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(4530))))  severity failure;
	assert RAM(4531) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(4531))))  severity failure;
	assert RAM(4532) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(4532))))  severity failure;
	assert RAM(4533) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(4533))))  severity failure;
	assert RAM(4534) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(4534))))  severity failure;
	assert RAM(4535) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(4535))))  severity failure;
	assert RAM(4536) = std_logic_vector(to_unsigned(72, 8)) report "TEST FALLITO (WORKING ZONE). Expected  72  found " & integer'image(to_integer(unsigned(RAM(4536))))  severity failure;
	assert RAM(4537) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(4537))))  severity failure;
	assert RAM(4538) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(4538))))  severity failure;
	assert RAM(4539) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(4539))))  severity failure;
	assert RAM(4540) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(4540))))  severity failure;
	assert RAM(4541) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(4541))))  severity failure;
	assert RAM(4542) = std_logic_vector(to_unsigned(185, 8)) report "TEST FALLITO (WORKING ZONE). Expected  185  found " & integer'image(to_integer(unsigned(RAM(4542))))  severity failure;
	assert RAM(4543) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(4543))))  severity failure;
	assert RAM(4544) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(4544))))  severity failure;
	assert RAM(4545) = std_logic_vector(to_unsigned(7, 8)) report "TEST FALLITO (WORKING ZONE). Expected  7  found " & integer'image(to_integer(unsigned(RAM(4545))))  severity failure;
	assert RAM(4546) = std_logic_vector(to_unsigned(24, 8)) report "TEST FALLITO (WORKING ZONE). Expected  24  found " & integer'image(to_integer(unsigned(RAM(4546))))  severity failure;
	assert RAM(4547) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(4547))))  severity failure;
	assert RAM(4548) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(4548))))  severity failure;
	assert RAM(4549) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(4549))))  severity failure;
	assert RAM(4550) = std_logic_vector(to_unsigned(182, 8)) report "TEST FALLITO (WORKING ZONE). Expected  182  found " & integer'image(to_integer(unsigned(RAM(4550))))  severity failure;
	assert RAM(4551) = std_logic_vector(to_unsigned(67, 8)) report "TEST FALLITO (WORKING ZONE). Expected  67  found " & integer'image(to_integer(unsigned(RAM(4551))))  severity failure;
	assert RAM(4552) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(4552))))  severity failure;
	assert RAM(4553) = std_logic_vector(to_unsigned(132, 8)) report "TEST FALLITO (WORKING ZONE). Expected  132  found " & integer'image(to_integer(unsigned(RAM(4553))))  severity failure;
	assert RAM(4554) = std_logic_vector(to_unsigned(147, 8)) report "TEST FALLITO (WORKING ZONE). Expected  147  found " & integer'image(to_integer(unsigned(RAM(4554))))  severity failure;
	assert RAM(4555) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(4555))))  severity failure;
	assert RAM(4556) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(4556))))  severity failure;
	assert RAM(4557) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(4557))))  severity failure;
	assert RAM(4558) = std_logic_vector(to_unsigned(105, 8)) report "TEST FALLITO (WORKING ZONE). Expected  105  found " & integer'image(to_integer(unsigned(RAM(4558))))  severity failure;
	assert RAM(4559) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(4559))))  severity failure;
	assert RAM(4560) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(4560))))  severity failure;
	assert RAM(4561) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(4561))))  severity failure;
	assert RAM(4562) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(4562))))  severity failure;
	assert RAM(4563) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(4563))))  severity failure;
	assert RAM(4564) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(4564))))  severity failure;
	assert RAM(4565) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(4565))))  severity failure;
	assert RAM(4566) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(4566))))  severity failure;
	assert RAM(4567) = std_logic_vector(to_unsigned(47, 8)) report "TEST FALLITO (WORKING ZONE). Expected  47  found " & integer'image(to_integer(unsigned(RAM(4567))))  severity failure;
	assert RAM(4568) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(4568))))  severity failure;
	assert RAM(4569) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(4569))))  severity failure;
	assert RAM(4570) = std_logic_vector(to_unsigned(203, 8)) report "TEST FALLITO (WORKING ZONE). Expected  203  found " & integer'image(to_integer(unsigned(RAM(4570))))  severity failure;
	assert RAM(4571) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(4571))))  severity failure;
	assert RAM(4572) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(4572))))  severity failure;
	assert RAM(4573) = std_logic_vector(to_unsigned(9, 8)) report "TEST FALLITO (WORKING ZONE). Expected  9  found " & integer'image(to_integer(unsigned(RAM(4573))))  severity failure;
	assert RAM(4574) = std_logic_vector(to_unsigned(225, 8)) report "TEST FALLITO (WORKING ZONE). Expected  225  found " & integer'image(to_integer(unsigned(RAM(4574))))  severity failure;
	assert RAM(4575) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(4575))))  severity failure;
	assert RAM(4576) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(4576))))  severity failure;
	assert RAM(4577) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(4577))))  severity failure;
	assert RAM(4578) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(4578))))  severity failure;
	assert RAM(4579) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(4579))))  severity failure;
	assert RAM(4580) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(4580))))  severity failure;
	assert RAM(4581) = std_logic_vector(to_unsigned(246, 8)) report "TEST FALLITO (WORKING ZONE). Expected  246  found " & integer'image(to_integer(unsigned(RAM(4581))))  severity failure;
	assert RAM(4582) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(4582))))  severity failure;
	assert RAM(4583) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(4583))))  severity failure;
	assert RAM(4584) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(4584))))  severity failure;
	assert RAM(4585) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(4585))))  severity failure;
	assert RAM(4586) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(4586))))  severity failure;
	assert RAM(4587) = std_logic_vector(to_unsigned(233, 8)) report "TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM(4587))))  severity failure;
	assert RAM(4588) = std_logic_vector(to_unsigned(25, 8)) report "TEST FALLITO (WORKING ZONE). Expected  25  found " & integer'image(to_integer(unsigned(RAM(4588))))  severity failure;
	assert RAM(4589) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(4589))))  severity failure;
	assert RAM(4590) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(4590))))  severity failure;
	assert RAM(4591) = std_logic_vector(to_unsigned(6, 8)) report "TEST FALLITO (WORKING ZONE). Expected  6  found " & integer'image(to_integer(unsigned(RAM(4591))))  severity failure;
	assert RAM(4592) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(4592))))  severity failure;
	assert RAM(4593) = std_logic_vector(to_unsigned(231, 8)) report "TEST FALLITO (WORKING ZONE). Expected  231  found " & integer'image(to_integer(unsigned(RAM(4593))))  severity failure;
	assert RAM(4594) = std_logic_vector(to_unsigned(234, 8)) report "TEST FALLITO (WORKING ZONE). Expected  234  found " & integer'image(to_integer(unsigned(RAM(4594))))  severity failure;
	assert RAM(4595) = std_logic_vector(to_unsigned(158, 8)) report "TEST FALLITO (WORKING ZONE). Expected  158  found " & integer'image(to_integer(unsigned(RAM(4595))))  severity failure;
	assert RAM(4596) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(4596))))  severity failure;
	assert RAM(4597) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(4597))))  severity failure;
	assert RAM(4598) = std_logic_vector(to_unsigned(254, 8)) report "TEST FALLITO (WORKING ZONE). Expected  254  found " & integer'image(to_integer(unsigned(RAM(4598))))  severity failure;
	assert RAM(4599) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(4599))))  severity failure;
	assert RAM(4600) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(4600))))  severity failure;
	assert RAM(4601) = std_logic_vector(to_unsigned(64, 8)) report "TEST FALLITO (WORKING ZONE). Expected  64  found " & integer'image(to_integer(unsigned(RAM(4601))))  severity failure;
	assert RAM(4602) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(4602))))  severity failure;
	assert RAM(4603) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(4603))))  severity failure;
	assert RAM(4604) = std_logic_vector(to_unsigned(42, 8)) report "TEST FALLITO (WORKING ZONE). Expected  42  found " & integer'image(to_integer(unsigned(RAM(4604))))  severity failure;
	assert RAM(4605) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(4605))))  severity failure;
	assert RAM(4606) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(4606))))  severity failure;
	assert RAM(4607) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(4607))))  severity failure;
	assert RAM(4608) = std_logic_vector(to_unsigned(136, 8)) report "TEST FALLITO (WORKING ZONE). Expected  136  found " & integer'image(to_integer(unsigned(RAM(4608))))  severity failure;
	assert RAM(4609) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(4609))))  severity failure;
	assert RAM(4610) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(4610))))  severity failure;
	assert RAM(4611) = std_logic_vector(to_unsigned(84, 8)) report "TEST FALLITO (WORKING ZONE). Expected  84  found " & integer'image(to_integer(unsigned(RAM(4611))))  severity failure;
	assert RAM(4612) = std_logic_vector(to_unsigned(226, 8)) report "TEST FALLITO (WORKING ZONE). Expected  226  found " & integer'image(to_integer(unsigned(RAM(4612))))  severity failure;
	assert RAM(4613) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(4613))))  severity failure;
	assert RAM(4614) = std_logic_vector(to_unsigned(81, 8)) report "TEST FALLITO (WORKING ZONE). Expected  81  found " & integer'image(to_integer(unsigned(RAM(4614))))  severity failure;
	assert RAM(4615) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(4615))))  severity failure;
	assert RAM(4616) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(4616))))  severity failure;
	assert RAM(4617) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(4617))))  severity failure;
	assert RAM(4618) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(4618))))  severity failure;
	assert RAM(4619) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(4619))))  severity failure;
	assert RAM(4620) = std_logic_vector(to_unsigned(133, 8)) report "TEST FALLITO (WORKING ZONE). Expected  133  found " & integer'image(to_integer(unsigned(RAM(4620))))  severity failure;
	assert RAM(4621) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(4621))))  severity failure;
	assert RAM(4622) = std_logic_vector(to_unsigned(172, 8)) report "TEST FALLITO (WORKING ZONE). Expected  172  found " & integer'image(to_integer(unsigned(RAM(4622))))  severity failure;
	assert RAM(4623) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(4623))))  severity failure;
	assert RAM(4624) = std_logic_vector(to_unsigned(165, 8)) report "TEST FALLITO (WORKING ZONE). Expected  165  found " & integer'image(to_integer(unsigned(RAM(4624))))  severity failure;
	assert RAM(4625) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(4625))))  severity failure;
	assert RAM(4626) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(4626))))  severity failure;
	assert RAM(4627) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(4627))))  severity failure;
	assert RAM(4628) = std_logic_vector(to_unsigned(170, 8)) report "TEST FALLITO (WORKING ZONE). Expected  170  found " & integer'image(to_integer(unsigned(RAM(4628))))  severity failure;
	assert RAM(4629) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(4629))))  severity failure;
	assert RAM(4630) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(4630))))  severity failure;
	assert RAM(4631) = std_logic_vector(to_unsigned(32, 8)) report "TEST FALLITO (WORKING ZONE). Expected  32  found " & integer'image(to_integer(unsigned(RAM(4631))))  severity failure;
	assert RAM(4632) = std_logic_vector(to_unsigned(71, 8)) report "TEST FALLITO (WORKING ZONE). Expected  71  found " & integer'image(to_integer(unsigned(RAM(4632))))  severity failure;
	assert RAM(4633) = std_logic_vector(to_unsigned(239, 8)) report "TEST FALLITO (WORKING ZONE). Expected  239  found " & integer'image(to_integer(unsigned(RAM(4633))))  severity failure;
	assert RAM(4634) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(4634))))  severity failure;
	assert RAM(4635) = std_logic_vector(to_unsigned(228, 8)) report "TEST FALLITO (WORKING ZONE). Expected  228  found " & integer'image(to_integer(unsigned(RAM(4635))))  severity failure;
	assert RAM(4636) = std_logic_vector(to_unsigned(115, 8)) report "TEST FALLITO (WORKING ZONE). Expected  115  found " & integer'image(to_integer(unsigned(RAM(4636))))  severity failure;
	assert RAM(4637) = std_logic_vector(to_unsigned(14, 8)) report "TEST FALLITO (WORKING ZONE). Expected  14  found " & integer'image(to_integer(unsigned(RAM(4637))))  severity failure;
	assert RAM(4638) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(4638))))  severity failure;
	assert RAM(4639) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(4639))))  severity failure;
	assert RAM(4640) = std_logic_vector(to_unsigned(80, 8)) report "TEST FALLITO (WORKING ZONE). Expected  80  found " & integer'image(to_integer(unsigned(RAM(4640))))  severity failure;
	assert RAM(4641) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(4641))))  severity failure;
	assert RAM(4642) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(4642))))  severity failure;
	assert RAM(4643) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(4643))))  severity failure;
	assert RAM(4644) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(4644))))  severity failure;
	assert RAM(4645) = std_logic_vector(to_unsigned(61, 8)) report "TEST FALLITO (WORKING ZONE). Expected  61  found " & integer'image(to_integer(unsigned(RAM(4645))))  severity failure;
	assert RAM(4646) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(4646))))  severity failure;
	assert RAM(4647) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(4647))))  severity failure;
	assert RAM(4648) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(4648))))  severity failure;
	assert RAM(4649) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(4649))))  severity failure;
	assert RAM(4650) = std_logic_vector(to_unsigned(135, 8)) report "TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM(4650))))  severity failure;
	assert RAM(4651) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(4651))))  severity failure;
	assert RAM(4652) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(4652))))  severity failure;
	assert RAM(4653) = std_logic_vector(to_unsigned(252, 8)) report "TEST FALLITO (WORKING ZONE). Expected  252  found " & integer'image(to_integer(unsigned(RAM(4653))))  severity failure;
	assert RAM(4654) = std_logic_vector(to_unsigned(245, 8)) report "TEST FALLITO (WORKING ZONE). Expected  245  found " & integer'image(to_integer(unsigned(RAM(4654))))  severity failure;
	assert RAM(4655) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(4655))))  severity failure;
	assert RAM(4656) = std_logic_vector(to_unsigned(164, 8)) report "TEST FALLITO (WORKING ZONE). Expected  164  found " & integer'image(to_integer(unsigned(RAM(4656))))  severity failure;
	assert RAM(4657) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(4657))))  severity failure;
	assert RAM(4658) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(4658))))  severity failure;
	assert RAM(4659) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(4659))))  severity failure;
	assert RAM(4660) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(4660))))  severity failure;
	assert RAM(4661) = std_logic_vector(to_unsigned(248, 8)) report "TEST FALLITO (WORKING ZONE). Expected  248  found " & integer'image(to_integer(unsigned(RAM(4661))))  severity failure;
	assert RAM(4662) = std_logic_vector(to_unsigned(118, 8)) report "TEST FALLITO (WORKING ZONE). Expected  118  found " & integer'image(to_integer(unsigned(RAM(4662))))  severity failure;
	assert RAM(4663) = std_logic_vector(to_unsigned(30, 8)) report "TEST FALLITO (WORKING ZONE). Expected  30  found " & integer'image(to_integer(unsigned(RAM(4663))))  severity failure;
	assert RAM(4664) = std_logic_vector(to_unsigned(94, 8)) report "TEST FALLITO (WORKING ZONE). Expected  94  found " & integer'image(to_integer(unsigned(RAM(4664))))  severity failure;
	assert RAM(4665) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(4665))))  severity failure;
	assert RAM(4666) = std_logic_vector(to_unsigned(193, 8)) report "TEST FALLITO (WORKING ZONE). Expected  193  found " & integer'image(to_integer(unsigned(RAM(4666))))  severity failure;
	assert RAM(4667) = std_logic_vector(to_unsigned(137, 8)) report "TEST FALLITO (WORKING ZONE). Expected  137  found " & integer'image(to_integer(unsigned(RAM(4667))))  severity failure;
	assert RAM(4668) = std_logic_vector(to_unsigned(208, 8)) report "TEST FALLITO (WORKING ZONE). Expected  208  found " & integer'image(to_integer(unsigned(RAM(4668))))  severity failure;
	assert RAM(4669) = std_logic_vector(to_unsigned(140, 8)) report "TEST FALLITO (WORKING ZONE). Expected  140  found " & integer'image(to_integer(unsigned(RAM(4669))))  severity failure;
	assert RAM(4670) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(4670))))  severity failure;
	assert RAM(4671) = std_logic_vector(to_unsigned(236, 8)) report "TEST FALLITO (WORKING ZONE). Expected  236  found " & integer'image(to_integer(unsigned(RAM(4671))))  severity failure;
	assert RAM(4672) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(4672))))  severity failure;
	assert RAM(4673) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(4673))))  severity failure;
	assert RAM(4674) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(4674))))  severity failure;
	assert RAM(4675) = std_logic_vector(to_unsigned(22, 8)) report "TEST FALLITO (WORKING ZONE). Expected  22  found " & integer'image(to_integer(unsigned(RAM(4675))))  severity failure;
	assert RAM(4676) = std_logic_vector(to_unsigned(128, 8)) report "TEST FALLITO (WORKING ZONE). Expected  128  found " & integer'image(to_integer(unsigned(RAM(4676))))  severity failure;
	assert RAM(4677) = std_logic_vector(to_unsigned(221, 8)) report "TEST FALLITO (WORKING ZONE). Expected  221  found " & integer'image(to_integer(unsigned(RAM(4677))))  severity failure;
	assert RAM(4678) = std_logic_vector(to_unsigned(66, 8)) report "TEST FALLITO (WORKING ZONE). Expected  66  found " & integer'image(to_integer(unsigned(RAM(4678))))  severity failure;
	assert RAM(4679) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(4679))))  severity failure;
	assert RAM(4680) = std_logic_vector(to_unsigned(106, 8)) report "TEST FALLITO (WORKING ZONE). Expected  106  found " & integer'image(to_integer(unsigned(RAM(4680))))  severity failure;
	assert RAM(4681) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(4681))))  severity failure;
	assert RAM(4682) = std_logic_vector(to_unsigned(232, 8)) report "TEST FALLITO (WORKING ZONE). Expected  232  found " & integer'image(to_integer(unsigned(RAM(4682))))  severity failure;
	assert RAM(4683) = std_logic_vector(to_unsigned(219, 8)) report "TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM(4683))))  severity failure;
	assert RAM(4684) = std_logic_vector(to_unsigned(198, 8)) report "TEST FALLITO (WORKING ZONE). Expected  198  found " & integer'image(to_integer(unsigned(RAM(4684))))  severity failure;
	assert RAM(4685) = std_logic_vector(to_unsigned(83, 8)) report "TEST FALLITO (WORKING ZONE). Expected  83  found " & integer'image(to_integer(unsigned(RAM(4685))))  severity failure;
	assert RAM(4686) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(4686))))  severity failure;
	assert RAM(4687) = std_logic_vector(to_unsigned(0, 8)) report "TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM(4687))))  severity failure;
	assert RAM(4688) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(4688))))  severity failure;
	assert RAM(4689) = std_logic_vector(to_unsigned(139, 8)) report "TEST FALLITO (WORKING ZONE). Expected  139  found " & integer'image(to_integer(unsigned(RAM(4689))))  severity failure;
	assert RAM(4690) = std_logic_vector(to_unsigned(124, 8)) report "TEST FALLITO (WORKING ZONE). Expected  124  found " & integer'image(to_integer(unsigned(RAM(4690))))  severity failure;
	assert RAM(4691) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(4691))))  severity failure;
	assert RAM(4692) = std_logic_vector(to_unsigned(154, 8)) report "TEST FALLITO (WORKING ZONE). Expected  154  found " & integer'image(to_integer(unsigned(RAM(4692))))  severity failure;
	assert RAM(4693) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(4693))))  severity failure;
	assert RAM(4694) = std_logic_vector(to_unsigned(26, 8)) report "TEST FALLITO (WORKING ZONE). Expected  26  found " & integer'image(to_integer(unsigned(RAM(4694))))  severity failure;
	assert RAM(4695) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(4695))))  severity failure;
	assert RAM(4696) = std_logic_vector(to_unsigned(216, 8)) report "TEST FALLITO (WORKING ZONE). Expected  216  found " & integer'image(to_integer(unsigned(RAM(4696))))  severity failure;
	assert RAM(4697) = std_logic_vector(to_unsigned(10, 8)) report "TEST FALLITO (WORKING ZONE). Expected  10  found " & integer'image(to_integer(unsigned(RAM(4697))))  severity failure;
	assert RAM(4698) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(4698))))  severity failure;
	assert RAM(4699) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(4699))))  severity failure;
	assert RAM(4700) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(4700))))  severity failure;
	assert RAM(4701) = std_logic_vector(to_unsigned(15, 8)) report "TEST FALLITO (WORKING ZONE). Expected  15  found " & integer'image(to_integer(unsigned(RAM(4701))))  severity failure;
	assert RAM(4702) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(4702))))  severity failure;
	assert RAM(4703) = std_logic_vector(to_unsigned(79, 8)) report "TEST FALLITO (WORKING ZONE). Expected  79  found " & integer'image(to_integer(unsigned(RAM(4703))))  severity failure;
	assert RAM(4704) = std_logic_vector(to_unsigned(53, 8)) report "TEST FALLITO (WORKING ZONE). Expected  53  found " & integer'image(to_integer(unsigned(RAM(4704))))  severity failure;
	assert RAM(4705) = std_logic_vector(to_unsigned(244, 8)) report "TEST FALLITO (WORKING ZONE). Expected  244  found " & integer'image(to_integer(unsigned(RAM(4705))))  severity failure;
	assert RAM(4706) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(4706))))  severity failure;
	assert RAM(4707) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(4707))))  severity failure;
	assert RAM(4708) = std_logic_vector(to_unsigned(113, 8)) report "TEST FALLITO (WORKING ZONE). Expected  113  found " & integer'image(to_integer(unsigned(RAM(4708))))  severity failure;
	assert RAM(4709) = std_logic_vector(to_unsigned(222, 8)) report "TEST FALLITO (WORKING ZONE). Expected  222  found " & integer'image(to_integer(unsigned(RAM(4709))))  severity failure;
	assert RAM(4710) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(4710))))  severity failure;
	assert RAM(4711) = std_logic_vector(to_unsigned(12, 8)) report "TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM(4711))))  severity failure;
	assert RAM(4712) = std_logic_vector(to_unsigned(159, 8)) report "TEST FALLITO (WORKING ZONE). Expected  159  found " & integer'image(to_integer(unsigned(RAM(4712))))  severity failure;
	assert RAM(4713) = std_logic_vector(to_unsigned(11, 8)) report "TEST FALLITO (WORKING ZONE). Expected  11  found " & integer'image(to_integer(unsigned(RAM(4713))))  severity failure;
	assert RAM(4714) = std_logic_vector(to_unsigned(4, 8)) report "TEST FALLITO (WORKING ZONE). Expected  4  found " & integer'image(to_integer(unsigned(RAM(4714))))  severity failure;
	assert RAM(4715) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(4715))))  severity failure;
	assert RAM(4716) = std_logic_vector(to_unsigned(108, 8)) report "TEST FALLITO (WORKING ZONE). Expected  108  found " & integer'image(to_integer(unsigned(RAM(4716))))  severity failure;
	assert RAM(4717) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(4717))))  severity failure;
	assert RAM(4718) = std_logic_vector(to_unsigned(3, 8)) report "TEST FALLITO (WORKING ZONE). Expected  3  found " & integer'image(to_integer(unsigned(RAM(4718))))  severity failure;
	assert RAM(4719) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(4719))))  severity failure;
	assert RAM(4720) = std_logic_vector(to_unsigned(54, 8)) report "TEST FALLITO (WORKING ZONE). Expected  54  found " & integer'image(to_integer(unsigned(RAM(4720))))  severity failure;
	assert RAM(4721) = std_logic_vector(to_unsigned(169, 8)) report "TEST FALLITO (WORKING ZONE). Expected  169  found " & integer'image(to_integer(unsigned(RAM(4721))))  severity failure;
	assert RAM(4722) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(4722))))  severity failure;
	assert RAM(4723) = std_logic_vector(to_unsigned(223, 8)) report "TEST FALLITO (WORKING ZONE). Expected  223  found " & integer'image(to_integer(unsigned(RAM(4723))))  severity failure;
	assert RAM(4724) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(4724))))  severity failure;
	assert RAM(4725) = std_logic_vector(to_unsigned(93, 8)) report "TEST FALLITO (WORKING ZONE). Expected  93  found " & integer'image(to_integer(unsigned(RAM(4725))))  severity failure;
	assert RAM(4726) = std_logic_vector(to_unsigned(142, 8)) report "TEST FALLITO (WORKING ZONE). Expected  142  found " & integer'image(to_integer(unsigned(RAM(4726))))  severity failure;
	assert RAM(4727) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(4727))))  severity failure;
	assert RAM(4728) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(4728))))  severity failure;
	assert RAM(4729) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(4729))))  severity failure;
	assert RAM(4730) = std_logic_vector(to_unsigned(160, 8)) report "TEST FALLITO (WORKING ZONE). Expected  160  found " & integer'image(to_integer(unsigned(RAM(4730))))  severity failure;
	assert RAM(4731) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(4731))))  severity failure;
	assert RAM(4732) = std_logic_vector(to_unsigned(200, 8)) report "TEST FALLITO (WORKING ZONE). Expected  200  found " & integer'image(to_integer(unsigned(RAM(4732))))  severity failure;
	assert RAM(4733) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(4733))))  severity failure;
	assert RAM(4734) = std_logic_vector(to_unsigned(242, 8)) report "TEST FALLITO (WORKING ZONE). Expected  242  found " & integer'image(to_integer(unsigned(RAM(4734))))  severity failure;
	assert RAM(4735) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(4735))))  severity failure;
	assert RAM(4736) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(4736))))  severity failure;
	assert RAM(4737) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(4737))))  severity failure;
	assert RAM(4738) = std_logic_vector(to_unsigned(255, 8)) report "TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM(4738))))  severity failure;
	assert RAM(4739) = std_logic_vector(to_unsigned(211, 8)) report "TEST FALLITO (WORKING ZONE). Expected  211  found " & integer'image(to_integer(unsigned(RAM(4739))))  severity failure;
	assert RAM(4740) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(4740))))  severity failure;
	assert RAM(4741) = std_logic_vector(to_unsigned(92, 8)) report "TEST FALLITO (WORKING ZONE). Expected  92  found " & integer'image(to_integer(unsigned(RAM(4741))))  severity failure;
	assert RAM(4742) = std_logic_vector(to_unsigned(120, 8)) report "TEST FALLITO (WORKING ZONE). Expected  120  found " & integer'image(to_integer(unsigned(RAM(4742))))  severity failure;
	assert RAM(4743) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(4743))))  severity failure;
	assert RAM(4744) = std_logic_vector(to_unsigned(27, 8)) report "TEST FALLITO (WORKING ZONE). Expected  27  found " & integer'image(to_integer(unsigned(RAM(4744))))  severity failure;
	assert RAM(4745) = std_logic_vector(to_unsigned(96, 8)) report "TEST FALLITO (WORKING ZONE). Expected  96  found " & integer'image(to_integer(unsigned(RAM(4745))))  severity failure;
	assert RAM(4746) = std_logic_vector(to_unsigned(46, 8)) report "TEST FALLITO (WORKING ZONE). Expected  46  found " & integer'image(to_integer(unsigned(RAM(4746))))  severity failure;
	assert RAM(4747) = std_logic_vector(to_unsigned(192, 8)) report "TEST FALLITO (WORKING ZONE). Expected  192  found " & integer'image(to_integer(unsigned(RAM(4747))))  severity failure;
	assert RAM(4748) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(4748))))  severity failure;
	assert RAM(4749) = std_logic_vector(to_unsigned(5, 8)) report "TEST FALLITO (WORKING ZONE). Expected  5  found " & integer'image(to_integer(unsigned(RAM(4749))))  severity failure;
	assert RAM(4750) = std_logic_vector(to_unsigned(227, 8)) report "TEST FALLITO (WORKING ZONE). Expected  227  found " & integer'image(to_integer(unsigned(RAM(4750))))  severity failure;
	assert RAM(4751) = std_logic_vector(to_unsigned(101, 8)) report "TEST FALLITO (WORKING ZONE). Expected  101  found " & integer'image(to_integer(unsigned(RAM(4751))))  severity failure;
	assert RAM(4752) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(4752))))  severity failure;
	assert RAM(4753) = std_logic_vector(to_unsigned(229, 8)) report "TEST FALLITO (WORKING ZONE). Expected  229  found " & integer'image(to_integer(unsigned(RAM(4753))))  severity failure;
	assert RAM(4754) = std_logic_vector(to_unsigned(2, 8)) report "TEST FALLITO (WORKING ZONE). Expected  2  found " & integer'image(to_integer(unsigned(RAM(4754))))  severity failure;
	assert RAM(4755) = std_logic_vector(to_unsigned(116, 8)) report "TEST FALLITO (WORKING ZONE). Expected  116  found " & integer'image(to_integer(unsigned(RAM(4755))))  severity failure;
	assert RAM(4756) = std_logic_vector(to_unsigned(152, 8)) report "TEST FALLITO (WORKING ZONE). Expected  152  found " & integer'image(to_integer(unsigned(RAM(4756))))  severity failure;
	assert RAM(4757) = std_logic_vector(to_unsigned(23, 8)) report "TEST FALLITO (WORKING ZONE). Expected  23  found " & integer'image(to_integer(unsigned(RAM(4757))))  severity failure;
	assert RAM(4758) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(4758))))  severity failure;
	assert RAM(4759) = std_logic_vector(to_unsigned(100, 8)) report "TEST FALLITO (WORKING ZONE). Expected  100  found " & integer'image(to_integer(unsigned(RAM(4759))))  severity failure;
	assert RAM(4760) = std_logic_vector(to_unsigned(201, 8)) report "TEST FALLITO (WORKING ZONE). Expected  201  found " & integer'image(to_integer(unsigned(RAM(4760))))  severity failure;
	assert RAM(4761) = std_logic_vector(to_unsigned(202, 8)) report "TEST FALLITO (WORKING ZONE). Expected  202  found " & integer'image(to_integer(unsigned(RAM(4761))))  severity failure;
	assert RAM(4762) = std_logic_vector(to_unsigned(58, 8)) report "TEST FALLITO (WORKING ZONE). Expected  58  found " & integer'image(to_integer(unsigned(RAM(4762))))  severity failure;
	assert RAM(4763) = std_logic_vector(to_unsigned(156, 8)) report "TEST FALLITO (WORKING ZONE). Expected  156  found " & integer'image(to_integer(unsigned(RAM(4763))))  severity failure;
	assert RAM(4764) = std_logic_vector(to_unsigned(33, 8)) report "TEST FALLITO (WORKING ZONE). Expected  33  found " & integer'image(to_integer(unsigned(RAM(4764))))  severity failure;
	assert RAM(4765) = std_logic_vector(to_unsigned(117, 8)) report "TEST FALLITO (WORKING ZONE). Expected  117  found " & integer'image(to_integer(unsigned(RAM(4765))))  severity failure;
	assert RAM(4766) = std_logic_vector(to_unsigned(18, 8)) report "TEST FALLITO (WORKING ZONE). Expected  18  found " & integer'image(to_integer(unsigned(RAM(4766))))  severity failure;
	assert RAM(4767) = std_logic_vector(to_unsigned(213, 8)) report "TEST FALLITO (WORKING ZONE). Expected  213  found " & integer'image(to_integer(unsigned(RAM(4767))))  severity failure;
	assert RAM(4768) = std_logic_vector(to_unsigned(68, 8)) report "TEST FALLITO (WORKING ZONE). Expected  68  found " & integer'image(to_integer(unsigned(RAM(4768))))  severity failure;
	assert RAM(4769) = std_logic_vector(to_unsigned(215, 8)) report "TEST FALLITO (WORKING ZONE). Expected  215  found " & integer'image(to_integer(unsigned(RAM(4769))))  severity failure;
	assert RAM(4770) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(4770))))  severity failure;
	assert RAM(4771) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(4771))))  severity failure;
	assert RAM(4772) = std_logic_vector(to_unsigned(175, 8)) report "TEST FALLITO (WORKING ZONE). Expected  175  found " & integer'image(to_integer(unsigned(RAM(4772))))  severity failure;
	assert RAM(4773) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(4773))))  severity failure;
	assert RAM(4774) = std_logic_vector(to_unsigned(1, 8)) report "TEST FALLITO (WORKING ZONE). Expected  1  found " & integer'image(to_integer(unsigned(RAM(4774))))  severity failure;
	assert RAM(4775) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(4775))))  severity failure;
	assert RAM(4776) = std_logic_vector(to_unsigned(161, 8)) report "TEST FALLITO (WORKING ZONE). Expected  161  found " & integer'image(to_integer(unsigned(RAM(4776))))  severity failure;
	assert RAM(4777) = std_logic_vector(to_unsigned(34, 8)) report "TEST FALLITO (WORKING ZONE). Expected  34  found " & integer'image(to_integer(unsigned(RAM(4777))))  severity failure;
	assert RAM(4778) = std_logic_vector(to_unsigned(123, 8)) report "TEST FALLITO (WORKING ZONE). Expected  123  found " & integer'image(to_integer(unsigned(RAM(4778))))  severity failure;
	assert RAM(4779) = std_logic_vector(to_unsigned(63, 8)) report "TEST FALLITO (WORKING ZONE). Expected  63  found " & integer'image(to_integer(unsigned(RAM(4779))))  severity failure;
	assert RAM(4780) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(4780))))  severity failure;
	assert RAM(4781) = std_logic_vector(to_unsigned(19, 8)) report "TEST FALLITO (WORKING ZONE). Expected  19  found " & integer'image(to_integer(unsigned(RAM(4781))))  severity failure;
	assert RAM(4782) = std_logic_vector(to_unsigned(163, 8)) report "TEST FALLITO (WORKING ZONE). Expected  163  found " & integer'image(to_integer(unsigned(RAM(4782))))  severity failure;
	assert RAM(4783) = std_logic_vector(to_unsigned(188, 8)) report "TEST FALLITO (WORKING ZONE). Expected  188  found " & integer'image(to_integer(unsigned(RAM(4783))))  severity failure;
	assert RAM(4784) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(4784))))  severity failure;
	assert RAM(4785) = std_logic_vector(to_unsigned(95, 8)) report "TEST FALLITO (WORKING ZONE). Expected  95  found " & integer'image(to_integer(unsigned(RAM(4785))))  severity failure;
	assert RAM(4786) = std_logic_vector(to_unsigned(74, 8)) report "TEST FALLITO (WORKING ZONE). Expected  74  found " & integer'image(to_integer(unsigned(RAM(4786))))  severity failure;
	assert RAM(4787) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(4787))))  severity failure;
	assert RAM(4788) = std_logic_vector(to_unsigned(52, 8)) report "TEST FALLITO (WORKING ZONE). Expected  52  found " & integer'image(to_integer(unsigned(RAM(4788))))  severity failure;
	assert RAM(4789) = std_logic_vector(to_unsigned(250, 8)) report "TEST FALLITO (WORKING ZONE). Expected  250  found " & integer'image(to_integer(unsigned(RAM(4789))))  severity failure;
	assert RAM(4790) = std_logic_vector(to_unsigned(109, 8)) report "TEST FALLITO (WORKING ZONE). Expected  109  found " & integer'image(to_integer(unsigned(RAM(4790))))  severity failure;
	assert RAM(4791) = std_logic_vector(to_unsigned(82, 8)) report "TEST FALLITO (WORKING ZONE). Expected  82  found " & integer'image(to_integer(unsigned(RAM(4791))))  severity failure;
	assert RAM(4792) = std_logic_vector(to_unsigned(48, 8)) report "TEST FALLITO (WORKING ZONE). Expected  48  found " & integer'image(to_integer(unsigned(RAM(4792))))  severity failure;
	assert RAM(4793) = std_logic_vector(to_unsigned(103, 8)) report "TEST FALLITO (WORKING ZONE). Expected  103  found " & integer'image(to_integer(unsigned(RAM(4793))))  severity failure;
	assert RAM(4794) = std_logic_vector(to_unsigned(179, 8)) report "TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM(4794))))  severity failure;
	assert RAM(4795) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(4795))))  severity failure;
	assert RAM(4796) = std_logic_vector(to_unsigned(217, 8)) report "TEST FALLITO (WORKING ZONE). Expected  217  found " & integer'image(to_integer(unsigned(RAM(4796))))  severity failure;
	assert RAM(4797) = std_logic_vector(to_unsigned(65, 8)) report "TEST FALLITO (WORKING ZONE). Expected  65  found " & integer'image(to_integer(unsigned(RAM(4797))))  severity failure;
	assert RAM(4798) = std_logic_vector(to_unsigned(247, 8)) report "TEST FALLITO (WORKING ZONE). Expected  247  found " & integer'image(to_integer(unsigned(RAM(4798))))  severity failure;
	assert RAM(4799) = std_logic_vector(to_unsigned(174, 8)) report "TEST FALLITO (WORKING ZONE). Expected  174  found " & integer'image(to_integer(unsigned(RAM(4799))))  severity failure;
	assert RAM(4800) = std_logic_vector(to_unsigned(189, 8)) report "TEST FALLITO (WORKING ZONE). Expected  189  found " & integer'image(to_integer(unsigned(RAM(4800))))  severity failure;
	assert RAM(4801) = std_logic_vector(to_unsigned(62, 8)) report "TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM(4801))))  severity failure;
	assert RAM(4802) = std_logic_vector(to_unsigned(122, 8)) report "TEST FALLITO (WORKING ZONE). Expected  122  found " & integer'image(to_integer(unsigned(RAM(4802))))  severity failure;
	assert RAM(4803) = std_logic_vector(to_unsigned(45, 8)) report "TEST FALLITO (WORKING ZONE). Expected  45  found " & integer'image(to_integer(unsigned(RAM(4803))))  severity failure;
	assert RAM(4804) = std_logic_vector(to_unsigned(238, 8)) report "TEST FALLITO (WORKING ZONE). Expected  238  found " & integer'image(to_integer(unsigned(RAM(4804))))  severity failure;
	assert RAM(4805) = std_logic_vector(to_unsigned(91, 8)) report "TEST FALLITO (WORKING ZONE). Expected  91  found " & integer'image(to_integer(unsigned(RAM(4805))))  severity failure;
	assert RAM(4806) = std_logic_vector(to_unsigned(177, 8)) report "TEST FALLITO (WORKING ZONE). Expected  177  found " & integer'image(to_integer(unsigned(RAM(4806))))  severity failure;
	assert RAM(4807) = std_logic_vector(to_unsigned(186, 8)) report "TEST FALLITO (WORKING ZONE). Expected  186  found " & integer'image(to_integer(unsigned(RAM(4807))))  severity failure;
	assert RAM(4808) = std_logic_vector(to_unsigned(240, 8)) report "TEST FALLITO (WORKING ZONE). Expected  240  found " & integer'image(to_integer(unsigned(RAM(4808))))  severity failure;
	assert RAM(4809) = std_logic_vector(to_unsigned(178, 8)) report "TEST FALLITO (WORKING ZONE). Expected  178  found " & integer'image(to_integer(unsigned(RAM(4809))))  severity failure;
	assert RAM(4810) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(4810))))  severity failure;
	assert RAM(4811) = std_logic_vector(to_unsigned(98, 8)) report "TEST FALLITO (WORKING ZONE). Expected  98  found " & integer'image(to_integer(unsigned(RAM(4811))))  severity failure;
	assert RAM(4812) = std_logic_vector(to_unsigned(153, 8)) report "TEST FALLITO (WORKING ZONE). Expected  153  found " & integer'image(to_integer(unsigned(RAM(4812))))  severity failure;
	assert RAM(4813) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(4813))))  severity failure;
	assert RAM(4814) = std_logic_vector(to_unsigned(251, 8)) report "TEST FALLITO (WORKING ZONE). Expected  251  found " & integer'image(to_integer(unsigned(RAM(4814))))  severity failure;
	assert RAM(4815) = std_logic_vector(to_unsigned(243, 8)) report "TEST FALLITO (WORKING ZONE). Expected  243  found " & integer'image(to_integer(unsigned(RAM(4815))))  severity failure;
	assert RAM(4816) = std_logic_vector(to_unsigned(76, 8)) report "TEST FALLITO (WORKING ZONE). Expected  76  found " & integer'image(to_integer(unsigned(RAM(4816))))  severity failure;
	assert RAM(4817) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(4817))))  severity failure;
	assert RAM(4818) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(4818))))  severity failure;
	assert RAM(4819) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(4819))))  severity failure;
	assert RAM(4820) = std_logic_vector(to_unsigned(56, 8)) report "TEST FALLITO (WORKING ZONE). Expected  56  found " & integer'image(to_integer(unsigned(RAM(4820))))  severity failure;
	assert RAM(4821) = std_logic_vector(to_unsigned(214, 8)) report "TEST FALLITO (WORKING ZONE). Expected  214  found " & integer'image(to_integer(unsigned(RAM(4821))))  severity failure;
	assert RAM(4822) = std_logic_vector(to_unsigned(111, 8)) report "TEST FALLITO (WORKING ZONE). Expected  111  found " & integer'image(to_integer(unsigned(RAM(4822))))  severity failure;
	assert RAM(4823) = std_logic_vector(to_unsigned(88, 8)) report "TEST FALLITO (WORKING ZONE). Expected  88  found " & integer'image(to_integer(unsigned(RAM(4823))))  severity failure;
	assert RAM(4824) = std_logic_vector(to_unsigned(50, 8)) report "TEST FALLITO (WORKING ZONE). Expected  50  found " & integer'image(to_integer(unsigned(RAM(4824))))  severity failure;
	assert RAM(4825) = std_logic_vector(to_unsigned(205, 8)) report "TEST FALLITO (WORKING ZONE). Expected  205  found " & integer'image(to_integer(unsigned(RAM(4825))))  severity failure;
	assert RAM(4826) = std_logic_vector(to_unsigned(146, 8)) report "TEST FALLITO (WORKING ZONE). Expected  146  found " & integer'image(to_integer(unsigned(RAM(4826))))  severity failure;
	assert RAM(4827) = std_logic_vector(to_unsigned(210, 8)) report "TEST FALLITO (WORKING ZONE). Expected  210  found " & integer'image(to_integer(unsigned(RAM(4827))))  severity failure;
	assert RAM(4828) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(4828))))  severity failure;
	assert RAM(4829) = std_logic_vector(to_unsigned(97, 8)) report "TEST FALLITO (WORKING ZONE). Expected  97  found " & integer'image(to_integer(unsigned(RAM(4829))))  severity failure;
	assert RAM(4830) = std_logic_vector(to_unsigned(197, 8)) report "TEST FALLITO (WORKING ZONE). Expected  197  found " & integer'image(to_integer(unsigned(RAM(4830))))  severity failure;
	assert RAM(4831) = std_logic_vector(to_unsigned(181, 8)) report "TEST FALLITO (WORKING ZONE). Expected  181  found " & integer'image(to_integer(unsigned(RAM(4831))))  severity failure;
	assert RAM(4832) = std_logic_vector(to_unsigned(167, 8)) report "TEST FALLITO (WORKING ZONE). Expected  167  found " & integer'image(to_integer(unsigned(RAM(4832))))  severity failure;
	assert RAM(4833) = std_logic_vector(to_unsigned(107, 8)) report "TEST FALLITO (WORKING ZONE). Expected  107  found " & integer'image(to_integer(unsigned(RAM(4833))))  severity failure;
	assert RAM(4834) = std_logic_vector(to_unsigned(114, 8)) report "TEST FALLITO (WORKING ZONE). Expected  114  found " & integer'image(to_integer(unsigned(RAM(4834))))  severity failure;
	assert RAM(4835) = std_logic_vector(to_unsigned(230, 8)) report "TEST FALLITO (WORKING ZONE). Expected  230  found " & integer'image(to_integer(unsigned(RAM(4835))))  severity failure;
	assert RAM(4836) = std_logic_vector(to_unsigned(44, 8)) report "TEST FALLITO (WORKING ZONE). Expected  44  found " & integer'image(to_integer(unsigned(RAM(4836))))  severity failure;
	assert RAM(4837) = std_logic_vector(to_unsigned(70, 8)) report "TEST FALLITO (WORKING ZONE). Expected  70  found " & integer'image(to_integer(unsigned(RAM(4837))))  severity failure;
	assert RAM(4838) = std_logic_vector(to_unsigned(190, 8)) report "TEST FALLITO (WORKING ZONE). Expected  190  found " & integer'image(to_integer(unsigned(RAM(4838))))  severity failure;
	assert RAM(4839) = std_logic_vector(to_unsigned(173, 8)) report "TEST FALLITO (WORKING ZONE). Expected  173  found " & integer'image(to_integer(unsigned(RAM(4839))))  severity failure;
	assert RAM(4840) = std_logic_vector(to_unsigned(180, 8)) report "TEST FALLITO (WORKING ZONE). Expected  180  found " & integer'image(to_integer(unsigned(RAM(4840))))  severity failure;
	assert RAM(4841) = std_logic_vector(to_unsigned(148, 8)) report "TEST FALLITO (WORKING ZONE). Expected  148  found " & integer'image(to_integer(unsigned(RAM(4841))))  severity failure;
	assert RAM(4842) = std_logic_vector(to_unsigned(130, 8)) report "TEST FALLITO (WORKING ZONE). Expected  130  found " & integer'image(to_integer(unsigned(RAM(4842))))  severity failure;
	assert RAM(4843) = std_logic_vector(to_unsigned(112, 8)) report "TEST FALLITO (WORKING ZONE). Expected  112  found " & integer'image(to_integer(unsigned(RAM(4843))))  severity failure;
	assert RAM(4844) = std_logic_vector(to_unsigned(90, 8)) report "TEST FALLITO (WORKING ZONE). Expected  90  found " & integer'image(to_integer(unsigned(RAM(4844))))  severity failure;
	assert RAM(4845) = std_logic_vector(to_unsigned(40, 8)) report "TEST FALLITO (WORKING ZONE). Expected  40  found " & integer'image(to_integer(unsigned(RAM(4845))))  severity failure;
	assert RAM(4846) = std_logic_vector(to_unsigned(36, 8)) report "TEST FALLITO (WORKING ZONE). Expected  36  found " & integer'image(to_integer(unsigned(RAM(4846))))  severity failure;
	assert RAM(4847) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(4847))))  severity failure;
	assert RAM(4848) = std_logic_vector(to_unsigned(55, 8)) report "TEST FALLITO (WORKING ZONE). Expected  55  found " & integer'image(to_integer(unsigned(RAM(4848))))  severity failure;
	assert RAM(4849) = std_logic_vector(to_unsigned(196, 8)) report "TEST FALLITO (WORKING ZONE). Expected  196  found " & integer'image(to_integer(unsigned(RAM(4849))))  severity failure;
	assert RAM(4850) = std_logic_vector(to_unsigned(166, 8)) report "TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM(4850))))  severity failure;
	assert RAM(4851) = std_logic_vector(to_unsigned(20, 8)) report "TEST FALLITO (WORKING ZONE). Expected  20  found " & integer'image(to_integer(unsigned(RAM(4851))))  severity failure;
	assert RAM(4852) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(4852))))  severity failure;
	assert RAM(4853) = std_logic_vector(to_unsigned(141, 8)) report "TEST FALLITO (WORKING ZONE). Expected  141  found " & integer'image(to_integer(unsigned(RAM(4853))))  severity failure;
	assert RAM(4854) = std_logic_vector(to_unsigned(21, 8)) report "TEST FALLITO (WORKING ZONE). Expected  21  found " & integer'image(to_integer(unsigned(RAM(4854))))  severity failure;
	assert RAM(4855) = std_logic_vector(to_unsigned(206, 8)) report "TEST FALLITO (WORKING ZONE). Expected  206  found " & integer'image(to_integer(unsigned(RAM(4855))))  severity failure;
	assert RAM(4856) = std_logic_vector(to_unsigned(28, 8)) report "TEST FALLITO (WORKING ZONE). Expected  28  found " & integer'image(to_integer(unsigned(RAM(4856))))  severity failure;
	assert RAM(4857) = std_logic_vector(to_unsigned(209, 8)) report "TEST FALLITO (WORKING ZONE). Expected  209  found " & integer'image(to_integer(unsigned(RAM(4857))))  severity failure;
	assert RAM(4858) = std_logic_vector(to_unsigned(184, 8)) report "TEST FALLITO (WORKING ZONE). Expected  184  found " & integer'image(to_integer(unsigned(RAM(4858))))  severity failure;
	assert RAM(4859) = std_logic_vector(to_unsigned(102, 8)) report "TEST FALLITO (WORKING ZONE). Expected  102  found " & integer'image(to_integer(unsigned(RAM(4859))))  severity failure;
	assert RAM(4860) = std_logic_vector(to_unsigned(191, 8)) report "TEST FALLITO (WORKING ZONE). Expected  191  found " & integer'image(to_integer(unsigned(RAM(4860))))  severity failure;
	assert RAM(4861) = std_logic_vector(to_unsigned(155, 8)) report "TEST FALLITO (WORKING ZONE). Expected  155  found " & integer'image(to_integer(unsigned(RAM(4861))))  severity failure;
    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;
end projecttb;
